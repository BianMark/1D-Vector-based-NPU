##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Sat Mar 22 07:34:55 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16_out
  CLASS BLOCK ;
  SIZE 730.0000 BY 130.0000 ;
  FOREIGN sram_w16_out 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 363.0500 0.0000 363.1500 0.5200 ;
    END
  END clk
  PIN D[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 46.8500 0.0000 46.9500 0.5200 ;
    END
  END D[159]
  PIN D[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 50.8500 0.0000 50.9500 0.5200 ;
    END
  END D[158]
  PIN D[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 54.8500 0.0000 54.9500 0.5200 ;
    END
  END D[157]
  PIN D[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 58.8500 0.0000 58.9500 0.5200 ;
    END
  END D[156]
  PIN D[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 62.8500 0.0000 62.9500 0.5200 ;
    END
  END D[155]
  PIN D[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 66.8500 0.0000 66.9500 0.5200 ;
    END
  END D[154]
  PIN D[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 70.8500 0.0000 70.9500 0.5200 ;
    END
  END D[153]
  PIN D[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 74.8500 0.0000 74.9500 0.5200 ;
    END
  END D[152]
  PIN D[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 78.8500 0.0000 78.9500 0.5200 ;
    END
  END D[151]
  PIN D[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 82.8500 0.0000 82.9500 0.5200 ;
    END
  END D[150]
  PIN D[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 86.8500 0.0000 86.9500 0.5200 ;
    END
  END D[149]
  PIN D[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 90.8500 0.0000 90.9500 0.5200 ;
    END
  END D[148]
  PIN D[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 94.8500 0.0000 94.9500 0.5200 ;
    END
  END D[147]
  PIN D[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 98.8500 0.0000 98.9500 0.5200 ;
    END
  END D[146]
  PIN D[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 102.8500 0.0000 102.9500 0.5200 ;
    END
  END D[145]
  PIN D[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 106.8500 0.0000 106.9500 0.5200 ;
    END
  END D[144]
  PIN D[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 110.8500 0.0000 110.9500 0.5200 ;
    END
  END D[143]
  PIN D[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 114.8500 0.0000 114.9500 0.5200 ;
    END
  END D[142]
  PIN D[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 118.8500 0.0000 118.9500 0.5200 ;
    END
  END D[141]
  PIN D[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 122.8500 0.0000 122.9500 0.5200 ;
    END
  END D[140]
  PIN D[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 126.8500 0.0000 126.9500 0.5200 ;
    END
  END D[139]
  PIN D[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 130.8500 0.0000 130.9500 0.5200 ;
    END
  END D[138]
  PIN D[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 134.8500 0.0000 134.9500 0.5200 ;
    END
  END D[137]
  PIN D[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 138.8500 0.0000 138.9500 0.5200 ;
    END
  END D[136]
  PIN D[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 142.8500 0.0000 142.9500 0.5200 ;
    END
  END D[135]
  PIN D[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 146.8500 0.0000 146.9500 0.5200 ;
    END
  END D[134]
  PIN D[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 150.8500 0.0000 150.9500 0.5200 ;
    END
  END D[133]
  PIN D[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 154.8500 0.0000 154.9500 0.5200 ;
    END
  END D[132]
  PIN D[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 158.8500 0.0000 158.9500 0.5200 ;
    END
  END D[131]
  PIN D[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 162.8500 0.0000 162.9500 0.5200 ;
    END
  END D[130]
  PIN D[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 166.8500 0.0000 166.9500 0.5200 ;
    END
  END D[129]
  PIN D[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 170.8500 0.0000 170.9500 0.5200 ;
    END
  END D[128]
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 174.8500 0.0000 174.9500 0.5200 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 178.8500 0.0000 178.9500 0.5200 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 182.8500 0.0000 182.9500 0.5200 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 186.8500 0.0000 186.9500 0.5200 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 190.8500 0.0000 190.9500 0.5200 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 194.8500 0.0000 194.9500 0.5200 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 198.8500 0.0000 198.9500 0.5200 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 202.8500 0.0000 202.9500 0.5200 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 206.8500 0.0000 206.9500 0.5200 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 210.8500 0.0000 210.9500 0.5200 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 214.8500 0.0000 214.9500 0.5200 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 218.8500 0.0000 218.9500 0.5200 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 222.8500 0.0000 222.9500 0.5200 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 226.8500 0.0000 226.9500 0.5200 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 230.8500 0.0000 230.9500 0.5200 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 234.8500 0.0000 234.9500 0.5200 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 238.8500 0.0000 238.9500 0.5200 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 242.8500 0.0000 242.9500 0.5200 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 246.8500 0.0000 246.9500 0.5200 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 250.8500 0.0000 250.9500 0.5200 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 254.8500 0.0000 254.9500 0.5200 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 258.8500 0.0000 258.9500 0.5200 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 262.8500 0.0000 262.9500 0.5200 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 266.8500 0.0000 266.9500 0.5200 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 270.8500 0.0000 270.9500 0.5200 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 274.8500 0.0000 274.9500 0.5200 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 278.8500 0.0000 278.9500 0.5200 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 282.8500 0.0000 282.9500 0.5200 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 286.8500 0.0000 286.9500 0.5200 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 290.8500 0.0000 290.9500 0.5200 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 294.8500 0.0000 294.9500 0.5200 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 298.8500 0.0000 298.9500 0.5200 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 302.8500 0.0000 302.9500 0.5200 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 306.8500 0.0000 306.9500 0.5200 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 310.8500 0.0000 310.9500 0.5200 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 314.8500 0.0000 314.9500 0.5200 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 318.8500 0.0000 318.9500 0.5200 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 322.8500 0.0000 322.9500 0.5200 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 326.8500 0.0000 326.9500 0.5200 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 330.8500 0.0000 330.9500 0.5200 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 334.8500 0.0000 334.9500 0.5200 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 338.8500 0.0000 338.9500 0.5200 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 342.8500 0.0000 342.9500 0.5200 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 346.8500 0.0000 346.9500 0.5200 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 350.8500 0.0000 350.9500 0.5200 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 354.8500 0.0000 354.9500 0.5200 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 358.8500 0.0000 358.9500 0.5200 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 362.8500 0.0000 362.9500 0.5200 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 366.8500 0.0000 366.9500 0.5200 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 370.8500 0.0000 370.9500 0.5200 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 374.8500 0.0000 374.9500 0.5200 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 378.8500 0.0000 378.9500 0.5200 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 382.8500 0.0000 382.9500 0.5200 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 386.8500 0.0000 386.9500 0.5200 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 390.8500 0.0000 390.9500 0.5200 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 394.8500 0.0000 394.9500 0.5200 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 398.8500 0.0000 398.9500 0.5200 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 402.8500 0.0000 402.9500 0.5200 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 406.8500 0.0000 406.9500 0.5200 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 410.8500 0.0000 410.9500 0.5200 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 414.8500 0.0000 414.9500 0.5200 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 418.8500 0.0000 418.9500 0.5200 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 422.8500 0.0000 422.9500 0.5200 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 426.8500 0.0000 426.9500 0.5200 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 430.8500 0.0000 430.9500 0.5200 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 434.8500 0.0000 434.9500 0.5200 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 438.8500 0.0000 438.9500 0.5200 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 442.8500 0.0000 442.9500 0.5200 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 446.8500 0.0000 446.9500 0.5200 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 450.8500 0.0000 450.9500 0.5200 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 454.8500 0.0000 454.9500 0.5200 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 458.8500 0.0000 458.9500 0.5200 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 462.8500 0.0000 462.9500 0.5200 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 466.8500 0.0000 466.9500 0.5200 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 470.8500 0.0000 470.9500 0.5200 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 474.8500 0.0000 474.9500 0.5200 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 478.8500 0.0000 478.9500 0.5200 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 482.8500 0.0000 482.9500 0.5200 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 486.8500 0.0000 486.9500 0.5200 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 490.8500 0.0000 490.9500 0.5200 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 494.8500 0.0000 494.9500 0.5200 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 498.8500 0.0000 498.9500 0.5200 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 502.8500 0.0000 502.9500 0.5200 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 506.8500 0.0000 506.9500 0.5200 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 510.8500 0.0000 510.9500 0.5200 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 514.8500 0.0000 514.9500 0.5200 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 518.8500 0.0000 518.9500 0.5200 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 522.8500 0.0000 522.9500 0.5200 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 526.8500 0.0000 526.9500 0.5200 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 530.8500 0.0000 530.9500 0.5200 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 534.8500 0.0000 534.9500 0.5200 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 538.8500 0.0000 538.9500 0.5200 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 542.8500 0.0000 542.9500 0.5200 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 546.8500 0.0000 546.9500 0.5200 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 550.8500 0.0000 550.9500 0.5200 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 554.8500 0.0000 554.9500 0.5200 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 558.8500 0.0000 558.9500 0.5200 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 562.8500 0.0000 562.9500 0.5200 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 566.8500 0.0000 566.9500 0.5200 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 570.8500 0.0000 570.9500 0.5200 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 574.8500 0.0000 574.9500 0.5200 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 578.8500 0.0000 578.9500 0.5200 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 582.8500 0.0000 582.9500 0.5200 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 586.8500 0.0000 586.9500 0.5200 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 590.8500 0.0000 590.9500 0.5200 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 594.8500 0.0000 594.9500 0.5200 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 598.8500 0.0000 598.9500 0.5200 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 602.8500 0.0000 602.9500 0.5200 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 606.8500 0.0000 606.9500 0.5200 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 610.8500 0.0000 610.9500 0.5200 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 614.8500 0.0000 614.9500 0.5200 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 618.8500 0.0000 618.9500 0.5200 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 622.8500 0.0000 622.9500 0.5200 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 626.8500 0.0000 626.9500 0.5200 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 630.8500 0.0000 630.9500 0.5200 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 634.8500 0.0000 634.9500 0.5200 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 638.8500 0.0000 638.9500 0.5200 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 642.8500 0.0000 642.9500 0.5200 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 646.8500 0.0000 646.9500 0.5200 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 650.8500 0.0000 650.9500 0.5200 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 654.8500 0.0000 654.9500 0.5200 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 658.8500 0.0000 658.9500 0.5200 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 662.8500 0.0000 662.9500 0.5200 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 666.8500 0.0000 666.9500 0.5200 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 670.8500 0.0000 670.9500 0.5200 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 674.8500 0.0000 674.9500 0.5200 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 678.8500 0.0000 678.9500 0.5200 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 682.8500 0.0000 682.9500 0.5200 ;
    END
  END D[0]
  PIN Q[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 46.8500 129.4800 46.9500 130.0000 ;
    END
  END Q[159]
  PIN Q[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 50.8500 129.4800 50.9500 130.0000 ;
    END
  END Q[158]
  PIN Q[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 54.8500 129.4800 54.9500 130.0000 ;
    END
  END Q[157]
  PIN Q[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 58.8500 129.4800 58.9500 130.0000 ;
    END
  END Q[156]
  PIN Q[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 62.8500 129.4800 62.9500 130.0000 ;
    END
  END Q[155]
  PIN Q[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 66.8500 129.4800 66.9500 130.0000 ;
    END
  END Q[154]
  PIN Q[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 70.8500 129.4800 70.9500 130.0000 ;
    END
  END Q[153]
  PIN Q[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 74.8500 129.4800 74.9500 130.0000 ;
    END
  END Q[152]
  PIN Q[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 78.8500 129.4800 78.9500 130.0000 ;
    END
  END Q[151]
  PIN Q[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 82.8500 129.4800 82.9500 130.0000 ;
    END
  END Q[150]
  PIN Q[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 86.8500 129.4800 86.9500 130.0000 ;
    END
  END Q[149]
  PIN Q[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 90.8500 129.4800 90.9500 130.0000 ;
    END
  END Q[148]
  PIN Q[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 94.8500 129.4800 94.9500 130.0000 ;
    END
  END Q[147]
  PIN Q[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 98.8500 129.4800 98.9500 130.0000 ;
    END
  END Q[146]
  PIN Q[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 102.8500 129.4800 102.9500 130.0000 ;
    END
  END Q[145]
  PIN Q[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 106.8500 129.4800 106.9500 130.0000 ;
    END
  END Q[144]
  PIN Q[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 110.8500 129.4800 110.9500 130.0000 ;
    END
  END Q[143]
  PIN Q[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 114.8500 129.4800 114.9500 130.0000 ;
    END
  END Q[142]
  PIN Q[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 118.8500 129.4800 118.9500 130.0000 ;
    END
  END Q[141]
  PIN Q[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 122.8500 129.4800 122.9500 130.0000 ;
    END
  END Q[140]
  PIN Q[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 126.8500 129.4800 126.9500 130.0000 ;
    END
  END Q[139]
  PIN Q[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 130.8500 129.4800 130.9500 130.0000 ;
    END
  END Q[138]
  PIN Q[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 134.8500 129.4800 134.9500 130.0000 ;
    END
  END Q[137]
  PIN Q[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 138.8500 129.4800 138.9500 130.0000 ;
    END
  END Q[136]
  PIN Q[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 142.8500 129.4800 142.9500 130.0000 ;
    END
  END Q[135]
  PIN Q[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 146.8500 129.4800 146.9500 130.0000 ;
    END
  END Q[134]
  PIN Q[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 150.8500 129.4800 150.9500 130.0000 ;
    END
  END Q[133]
  PIN Q[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 154.8500 129.4800 154.9500 130.0000 ;
    END
  END Q[132]
  PIN Q[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 158.8500 129.4800 158.9500 130.0000 ;
    END
  END Q[131]
  PIN Q[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 162.8500 129.4800 162.9500 130.0000 ;
    END
  END Q[130]
  PIN Q[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 166.8500 129.4800 166.9500 130.0000 ;
    END
  END Q[129]
  PIN Q[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 170.8500 129.4800 170.9500 130.0000 ;
    END
  END Q[128]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 174.8500 129.4800 174.9500 130.0000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 178.8500 129.4800 178.9500 130.0000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 182.8500 129.4800 182.9500 130.0000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 186.8500 129.4800 186.9500 130.0000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 190.8500 129.4800 190.9500 130.0000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 194.8500 129.4800 194.9500 130.0000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 198.8500 129.4800 198.9500 130.0000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 202.8500 129.4800 202.9500 130.0000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 206.8500 129.4800 206.9500 130.0000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 210.8500 129.4800 210.9500 130.0000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 214.8500 129.4800 214.9500 130.0000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 218.8500 129.4800 218.9500 130.0000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 222.8500 129.4800 222.9500 130.0000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 226.8500 129.4800 226.9500 130.0000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 230.8500 129.4800 230.9500 130.0000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 234.8500 129.4800 234.9500 130.0000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 238.8500 129.4800 238.9500 130.0000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 242.8500 129.4800 242.9500 130.0000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 246.8500 129.4800 246.9500 130.0000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 250.8500 129.4800 250.9500 130.0000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 254.8500 129.4800 254.9500 130.0000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 258.8500 129.4800 258.9500 130.0000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 262.8500 129.4800 262.9500 130.0000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 266.8500 129.4800 266.9500 130.0000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 270.8500 129.4800 270.9500 130.0000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 274.8500 129.4800 274.9500 130.0000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 278.8500 129.4800 278.9500 130.0000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 282.8500 129.4800 282.9500 130.0000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 286.8500 129.4800 286.9500 130.0000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 290.8500 129.4800 290.9500 130.0000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 294.8500 129.4800 294.9500 130.0000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 298.8500 129.4800 298.9500 130.0000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 302.8500 129.4800 302.9500 130.0000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 306.8500 129.4800 306.9500 130.0000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 310.8500 129.4800 310.9500 130.0000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 314.8500 129.4800 314.9500 130.0000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 318.8500 129.4800 318.9500 130.0000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 322.8500 129.4800 322.9500 130.0000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 326.8500 129.4800 326.9500 130.0000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 330.8500 129.4800 330.9500 130.0000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 334.8500 129.4800 334.9500 130.0000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 338.8500 129.4800 338.9500 130.0000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 342.8500 129.4800 342.9500 130.0000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 346.8500 129.4800 346.9500 130.0000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 350.8500 129.4800 350.9500 130.0000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 354.8500 129.4800 354.9500 130.0000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 358.8500 129.4800 358.9500 130.0000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 362.8500 129.4800 362.9500 130.0000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 366.8500 129.4800 366.9500 130.0000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 370.8500 129.4800 370.9500 130.0000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 374.8500 129.4800 374.9500 130.0000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 378.8500 129.4800 378.9500 130.0000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 382.8500 129.4800 382.9500 130.0000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 386.8500 129.4800 386.9500 130.0000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 390.8500 129.4800 390.9500 130.0000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 394.8500 129.4800 394.9500 130.0000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 398.8500 129.4800 398.9500 130.0000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 402.8500 129.4800 402.9500 130.0000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 406.8500 129.4800 406.9500 130.0000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 410.8500 129.4800 410.9500 130.0000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 414.8500 129.4800 414.9500 130.0000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 418.8500 129.4800 418.9500 130.0000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 422.8500 129.4800 422.9500 130.0000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 426.8500 129.4800 426.9500 130.0000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 430.8500 129.4800 430.9500 130.0000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 434.8500 129.4800 434.9500 130.0000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 438.8500 129.4800 438.9500 130.0000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 442.8500 129.4800 442.9500 130.0000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 446.8500 129.4800 446.9500 130.0000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 450.8500 129.4800 450.9500 130.0000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 454.8500 129.4800 454.9500 130.0000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 458.8500 129.4800 458.9500 130.0000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 462.8500 129.4800 462.9500 130.0000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 466.8500 129.4800 466.9500 130.0000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 470.8500 129.4800 470.9500 130.0000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 474.8500 129.4800 474.9500 130.0000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 478.8500 129.4800 478.9500 130.0000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 482.8500 129.4800 482.9500 130.0000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 486.8500 129.4800 486.9500 130.0000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 490.8500 129.4800 490.9500 130.0000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 494.8500 129.4800 494.9500 130.0000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 498.8500 129.4800 498.9500 130.0000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 502.8500 129.4800 502.9500 130.0000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 506.8500 129.4800 506.9500 130.0000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 510.8500 129.4800 510.9500 130.0000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 514.8500 129.4800 514.9500 130.0000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 518.8500 129.4800 518.9500 130.0000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 522.8500 129.4800 522.9500 130.0000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 526.8500 129.4800 526.9500 130.0000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 530.8500 129.4800 530.9500 130.0000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 534.8500 129.4800 534.9500 130.0000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 538.8500 129.4800 538.9500 130.0000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 542.8500 129.4800 542.9500 130.0000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 546.8500 129.4800 546.9500 130.0000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 550.8500 129.4800 550.9500 130.0000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 554.8500 129.4800 554.9500 130.0000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 558.8500 129.4800 558.9500 130.0000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 562.8500 129.4800 562.9500 130.0000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 566.8500 129.4800 566.9500 130.0000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 570.8500 129.4800 570.9500 130.0000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 574.8500 129.4800 574.9500 130.0000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 578.8500 129.4800 578.9500 130.0000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 582.8500 129.4800 582.9500 130.0000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 586.8500 129.4800 586.9500 130.0000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 590.8500 129.4800 590.9500 130.0000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 594.8500 129.4800 594.9500 130.0000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 598.8500 129.4800 598.9500 130.0000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 602.8500 129.4800 602.9500 130.0000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 606.8500 129.4800 606.9500 130.0000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 610.8500 129.4800 610.9500 130.0000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 614.8500 129.4800 614.9500 130.0000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 618.8500 129.4800 618.9500 130.0000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 622.8500 129.4800 622.9500 130.0000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 626.8500 129.4800 626.9500 130.0000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 630.8500 129.4800 630.9500 130.0000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 634.8500 129.4800 634.9500 130.0000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 638.8500 129.4800 638.9500 130.0000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 642.8500 129.4800 642.9500 130.0000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 646.8500 129.4800 646.9500 130.0000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 650.8500 129.4800 650.9500 130.0000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 654.8500 129.4800 654.9500 130.0000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 658.8500 129.4800 658.9500 130.0000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 662.8500 129.4800 662.9500 130.0000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 666.8500 129.4800 666.9500 130.0000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 670.8500 129.4800 670.9500 130.0000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 674.8500 129.4800 674.9500 130.0000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 678.8500 129.4800 678.9500 130.0000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 682.8500 129.4800 682.9500 130.0000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 59.1500 0.5200 59.2500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 55.1500 0.5200 55.2500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 75.1500 0.5200 75.2500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 71.1500 0.5200 71.2500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 67.1500 0.5200 67.2500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 63.1500 0.5200 63.2500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 25.0000 15.0000 26.0000 115.0000 ;
        RECT 42.2300 15.0000 43.2300 115.0000 ;
        RECT 59.4600 15.0000 60.4600 115.0000 ;
        RECT 76.6900 15.0000 77.6900 115.0000 ;
        RECT 93.9200 15.0000 94.9200 115.0000 ;
        RECT 111.1500 15.0000 112.1500 115.0000 ;
        RECT 128.3800 15.0000 129.3800 115.0000 ;
        RECT 145.6100 15.0000 146.6100 115.0000 ;
        RECT 162.8400 15.0000 163.8400 115.0000 ;
        RECT 180.0700 15.0000 181.0700 115.0000 ;
        RECT 197.3000 15.0000 198.3000 115.0000 ;
        RECT 214.5300 15.0000 215.5300 115.0000 ;
        RECT 231.7600 15.0000 232.7600 115.0000 ;
        RECT 248.9900 15.0000 249.9900 115.0000 ;
        RECT 266.2200 15.0000 267.2200 115.0000 ;
        RECT 283.4500 15.0000 284.4500 115.0000 ;
        RECT 300.6800 15.0000 301.6800 115.0000 ;
        RECT 317.9100 15.0000 318.9100 115.0000 ;
        RECT 335.1400 15.0000 336.1400 115.0000 ;
        RECT 352.3700 15.0000 353.3700 115.0000 ;
        RECT 369.6000 15.0000 370.6000 115.0000 ;
        RECT 386.8300 15.0000 387.8300 115.0000 ;
        RECT 404.0600 15.0000 405.0600 115.0000 ;
        RECT 421.2900 15.0000 422.2900 115.0000 ;
        RECT 438.5200 15.0000 439.5200 115.0000 ;
        RECT 455.7500 15.0000 456.7500 115.0000 ;
        RECT 472.9800 15.0000 473.9800 115.0000 ;
        RECT 490.2100 15.0000 491.2100 115.0000 ;
        RECT 507.4400 15.0000 508.4400 115.0000 ;
        RECT 524.6700 15.0000 525.6700 115.0000 ;
        RECT 541.9000 15.0000 542.9000 115.0000 ;
        RECT 696.9700 15.0000 697.9700 115.0000 ;
        RECT 679.7400 15.0000 680.7400 115.0000 ;
        RECT 662.5100 15.0000 663.5100 115.0000 ;
        RECT 645.2800 15.0000 646.2800 115.0000 ;
        RECT 628.0500 15.0000 629.0500 115.0000 ;
        RECT 610.8200 15.0000 611.8200 115.0000 ;
        RECT 593.5900 15.0000 594.5900 115.0000 ;
        RECT 576.3600 15.0000 577.3600 115.0000 ;
        RECT 559.1300 15.0000 560.1300 115.0000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 182.0700 15.0000 183.0700 115.0000 ;
        RECT 164.8400 15.0000 165.8400 115.0000 ;
        RECT 147.6100 15.0000 148.6100 115.0000 ;
        RECT 130.3800 15.0000 131.3800 115.0000 ;
        RECT 113.1500 15.0000 114.1500 115.0000 ;
        RECT 95.9200 15.0000 96.9200 115.0000 ;
        RECT 78.6900 15.0000 79.6900 115.0000 ;
        RECT 61.4600 15.0000 62.4600 115.0000 ;
        RECT 44.2300 15.0000 45.2300 115.0000 ;
        RECT 27.0000 15.0000 28.0000 115.0000 ;
        RECT 199.3000 15.0000 200.3000 115.0000 ;
        RECT 216.5300 15.0000 217.5300 115.0000 ;
        RECT 233.7600 15.0000 234.7600 115.0000 ;
        RECT 250.9900 15.0000 251.9900 115.0000 ;
        RECT 268.2200 15.0000 269.2200 115.0000 ;
        RECT 285.4500 15.0000 286.4500 115.0000 ;
        RECT 302.6800 15.0000 303.6800 115.0000 ;
        RECT 319.9100 15.0000 320.9100 115.0000 ;
        RECT 337.1400 15.0000 338.1400 115.0000 ;
        RECT 354.3700 15.0000 355.3700 115.0000 ;
        RECT 526.6700 15.0000 527.6700 115.0000 ;
        RECT 509.4400 15.0000 510.4400 115.0000 ;
        RECT 492.2100 15.0000 493.2100 115.0000 ;
        RECT 474.9800 15.0000 475.9800 115.0000 ;
        RECT 457.7500 15.0000 458.7500 115.0000 ;
        RECT 440.5200 15.0000 441.5200 115.0000 ;
        RECT 423.2900 15.0000 424.2900 115.0000 ;
        RECT 406.0600 15.0000 407.0600 115.0000 ;
        RECT 388.8300 15.0000 389.8300 115.0000 ;
        RECT 371.6000 15.0000 372.6000 115.0000 ;
        RECT 543.9000 15.0000 544.9000 115.0000 ;
        RECT 561.1300 15.0000 562.1300 115.0000 ;
        RECT 578.3600 15.0000 579.3600 115.0000 ;
        RECT 595.5900 15.0000 596.5900 115.0000 ;
        RECT 612.8200 15.0000 613.8200 115.0000 ;
        RECT 630.0500 15.0000 631.0500 115.0000 ;
        RECT 647.2800 15.0000 648.2800 115.0000 ;
        RECT 664.5100 15.0000 665.5100 115.0000 ;
        RECT 681.7400 15.0000 682.7400 115.0000 ;
        RECT 698.9700 15.0000 699.9700 115.0000 ;
        RECT 182.0700 14.8350 183.0700 15.1650 ;
        RECT 27.0000 14.8350 28.0000 15.1650 ;
        RECT 44.2300 14.8350 45.2300 15.1650 ;
        RECT 61.4600 14.8350 62.4600 15.1650 ;
        RECT 78.6900 14.8350 79.6900 15.1650 ;
        RECT 113.1500 14.8350 114.1500 15.1650 ;
        RECT 95.9200 14.8350 96.9200 15.1650 ;
        RECT 130.3800 14.8350 131.3800 15.1650 ;
        RECT 147.6100 14.8350 148.6100 15.1650 ;
        RECT 164.8400 14.8350 165.8400 15.1650 ;
        RECT 199.3000 14.8350 200.3000 15.1650 ;
        RECT 216.5300 14.8350 217.5300 15.1650 ;
        RECT 233.7600 14.8350 234.7600 15.1650 ;
        RECT 268.2200 14.8350 269.2200 15.1650 ;
        RECT 250.9900 14.8350 251.9900 15.1650 ;
        RECT 285.4500 14.8350 286.4500 15.1650 ;
        RECT 302.6800 14.8350 303.6800 15.1650 ;
        RECT 337.1400 14.8350 338.1400 15.1650 ;
        RECT 319.9100 14.8350 320.9100 15.1650 ;
        RECT 354.3700 14.8350 355.3700 15.1650 ;
        RECT 371.6000 14.8350 372.6000 15.1650 ;
        RECT 406.0600 14.8350 407.0600 15.1650 ;
        RECT 388.8300 14.8350 389.8300 15.1650 ;
        RECT 423.2900 14.8350 424.2900 15.1650 ;
        RECT 440.5200 14.8350 441.5200 15.1650 ;
        RECT 474.9800 14.8350 475.9800 15.1650 ;
        RECT 457.7500 14.8350 458.7500 15.1650 ;
        RECT 492.2100 14.8350 493.2100 15.1650 ;
        RECT 509.4400 14.8350 510.4400 15.1650 ;
        RECT 543.9000 14.8350 544.9000 15.1650 ;
        RECT 526.6700 14.8350 527.6700 15.1650 ;
        RECT 561.1300 14.8350 562.1300 15.1650 ;
        RECT 578.3600 14.8350 579.3600 15.1650 ;
        RECT 595.5900 14.8350 596.5900 15.1650 ;
        RECT 612.8200 14.8350 613.8200 15.1650 ;
        RECT 630.0500 14.8350 631.0500 15.1650 ;
        RECT 647.2800 14.8350 648.2800 15.1650 ;
        RECT 664.5100 14.8350 665.5100 15.1650 ;
        RECT 681.7400 14.8350 682.7400 15.1650 ;
        RECT 698.9700 14.8350 699.9700 15.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 730.0000 130.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.6200 730.0000 130.0000 ;
      RECT 363.2500 0.0000 730.0000 0.6200 ;
      RECT 0.0000 0.0000 362.9500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 75.3500 730.0000 130.0000 ;
      RECT 0.6200 75.0500 730.0000 75.3500 ;
      RECT 0.0000 71.3500 730.0000 75.0500 ;
      RECT 0.6200 71.0500 730.0000 71.3500 ;
      RECT 0.0000 67.3500 730.0000 71.0500 ;
      RECT 0.6200 67.0500 730.0000 67.3500 ;
      RECT 0.0000 63.3500 730.0000 67.0500 ;
      RECT 0.6200 63.0500 730.0000 63.3500 ;
      RECT 0.0000 59.3500 730.0000 63.0500 ;
      RECT 0.6200 59.0500 730.0000 59.3500 ;
      RECT 0.0000 55.3500 730.0000 59.0500 ;
      RECT 0.6200 55.0500 730.0000 55.3500 ;
      RECT 0.0000 0.0000 730.0000 55.0500 ;
    LAYER M4 ;
      RECT 683.0500 129.3800 730.0000 130.0000 ;
      RECT 679.0500 129.3800 682.7500 130.0000 ;
      RECT 675.0500 129.3800 678.7500 130.0000 ;
      RECT 671.0500 129.3800 674.7500 130.0000 ;
      RECT 667.0500 129.3800 670.7500 130.0000 ;
      RECT 663.0500 129.3800 666.7500 130.0000 ;
      RECT 659.0500 129.3800 662.7500 130.0000 ;
      RECT 655.0500 129.3800 658.7500 130.0000 ;
      RECT 651.0500 129.3800 654.7500 130.0000 ;
      RECT 647.0500 129.3800 650.7500 130.0000 ;
      RECT 643.0500 129.3800 646.7500 130.0000 ;
      RECT 639.0500 129.3800 642.7500 130.0000 ;
      RECT 635.0500 129.3800 638.7500 130.0000 ;
      RECT 631.0500 129.3800 634.7500 130.0000 ;
      RECT 627.0500 129.3800 630.7500 130.0000 ;
      RECT 623.0500 129.3800 626.7500 130.0000 ;
      RECT 619.0500 129.3800 622.7500 130.0000 ;
      RECT 615.0500 129.3800 618.7500 130.0000 ;
      RECT 611.0500 129.3800 614.7500 130.0000 ;
      RECT 607.0500 129.3800 610.7500 130.0000 ;
      RECT 603.0500 129.3800 606.7500 130.0000 ;
      RECT 599.0500 129.3800 602.7500 130.0000 ;
      RECT 595.0500 129.3800 598.7500 130.0000 ;
      RECT 591.0500 129.3800 594.7500 130.0000 ;
      RECT 587.0500 129.3800 590.7500 130.0000 ;
      RECT 583.0500 129.3800 586.7500 130.0000 ;
      RECT 579.0500 129.3800 582.7500 130.0000 ;
      RECT 575.0500 129.3800 578.7500 130.0000 ;
      RECT 571.0500 129.3800 574.7500 130.0000 ;
      RECT 567.0500 129.3800 570.7500 130.0000 ;
      RECT 563.0500 129.3800 566.7500 130.0000 ;
      RECT 559.0500 129.3800 562.7500 130.0000 ;
      RECT 555.0500 129.3800 558.7500 130.0000 ;
      RECT 551.0500 129.3800 554.7500 130.0000 ;
      RECT 547.0500 129.3800 550.7500 130.0000 ;
      RECT 543.0500 129.3800 546.7500 130.0000 ;
      RECT 539.0500 129.3800 542.7500 130.0000 ;
      RECT 535.0500 129.3800 538.7500 130.0000 ;
      RECT 531.0500 129.3800 534.7500 130.0000 ;
      RECT 527.0500 129.3800 530.7500 130.0000 ;
      RECT 523.0500 129.3800 526.7500 130.0000 ;
      RECT 519.0500 129.3800 522.7500 130.0000 ;
      RECT 515.0500 129.3800 518.7500 130.0000 ;
      RECT 511.0500 129.3800 514.7500 130.0000 ;
      RECT 507.0500 129.3800 510.7500 130.0000 ;
      RECT 503.0500 129.3800 506.7500 130.0000 ;
      RECT 499.0500 129.3800 502.7500 130.0000 ;
      RECT 495.0500 129.3800 498.7500 130.0000 ;
      RECT 491.0500 129.3800 494.7500 130.0000 ;
      RECT 487.0500 129.3800 490.7500 130.0000 ;
      RECT 483.0500 129.3800 486.7500 130.0000 ;
      RECT 479.0500 129.3800 482.7500 130.0000 ;
      RECT 475.0500 129.3800 478.7500 130.0000 ;
      RECT 471.0500 129.3800 474.7500 130.0000 ;
      RECT 467.0500 129.3800 470.7500 130.0000 ;
      RECT 463.0500 129.3800 466.7500 130.0000 ;
      RECT 459.0500 129.3800 462.7500 130.0000 ;
      RECT 455.0500 129.3800 458.7500 130.0000 ;
      RECT 451.0500 129.3800 454.7500 130.0000 ;
      RECT 447.0500 129.3800 450.7500 130.0000 ;
      RECT 443.0500 129.3800 446.7500 130.0000 ;
      RECT 439.0500 129.3800 442.7500 130.0000 ;
      RECT 435.0500 129.3800 438.7500 130.0000 ;
      RECT 431.0500 129.3800 434.7500 130.0000 ;
      RECT 427.0500 129.3800 430.7500 130.0000 ;
      RECT 423.0500 129.3800 426.7500 130.0000 ;
      RECT 419.0500 129.3800 422.7500 130.0000 ;
      RECT 415.0500 129.3800 418.7500 130.0000 ;
      RECT 411.0500 129.3800 414.7500 130.0000 ;
      RECT 407.0500 129.3800 410.7500 130.0000 ;
      RECT 403.0500 129.3800 406.7500 130.0000 ;
      RECT 399.0500 129.3800 402.7500 130.0000 ;
      RECT 395.0500 129.3800 398.7500 130.0000 ;
      RECT 391.0500 129.3800 394.7500 130.0000 ;
      RECT 387.0500 129.3800 390.7500 130.0000 ;
      RECT 383.0500 129.3800 386.7500 130.0000 ;
      RECT 379.0500 129.3800 382.7500 130.0000 ;
      RECT 375.0500 129.3800 378.7500 130.0000 ;
      RECT 371.0500 129.3800 374.7500 130.0000 ;
      RECT 367.0500 129.3800 370.7500 130.0000 ;
      RECT 363.0500 129.3800 366.7500 130.0000 ;
      RECT 359.0500 129.3800 362.7500 130.0000 ;
      RECT 355.0500 129.3800 358.7500 130.0000 ;
      RECT 351.0500 129.3800 354.7500 130.0000 ;
      RECT 347.0500 129.3800 350.7500 130.0000 ;
      RECT 343.0500 129.3800 346.7500 130.0000 ;
      RECT 339.0500 129.3800 342.7500 130.0000 ;
      RECT 335.0500 129.3800 338.7500 130.0000 ;
      RECT 331.0500 129.3800 334.7500 130.0000 ;
      RECT 327.0500 129.3800 330.7500 130.0000 ;
      RECT 323.0500 129.3800 326.7500 130.0000 ;
      RECT 319.0500 129.3800 322.7500 130.0000 ;
      RECT 315.0500 129.3800 318.7500 130.0000 ;
      RECT 311.0500 129.3800 314.7500 130.0000 ;
      RECT 307.0500 129.3800 310.7500 130.0000 ;
      RECT 303.0500 129.3800 306.7500 130.0000 ;
      RECT 299.0500 129.3800 302.7500 130.0000 ;
      RECT 295.0500 129.3800 298.7500 130.0000 ;
      RECT 291.0500 129.3800 294.7500 130.0000 ;
      RECT 287.0500 129.3800 290.7500 130.0000 ;
      RECT 283.0500 129.3800 286.7500 130.0000 ;
      RECT 279.0500 129.3800 282.7500 130.0000 ;
      RECT 275.0500 129.3800 278.7500 130.0000 ;
      RECT 271.0500 129.3800 274.7500 130.0000 ;
      RECT 267.0500 129.3800 270.7500 130.0000 ;
      RECT 263.0500 129.3800 266.7500 130.0000 ;
      RECT 259.0500 129.3800 262.7500 130.0000 ;
      RECT 255.0500 129.3800 258.7500 130.0000 ;
      RECT 251.0500 129.3800 254.7500 130.0000 ;
      RECT 247.0500 129.3800 250.7500 130.0000 ;
      RECT 243.0500 129.3800 246.7500 130.0000 ;
      RECT 239.0500 129.3800 242.7500 130.0000 ;
      RECT 235.0500 129.3800 238.7500 130.0000 ;
      RECT 231.0500 129.3800 234.7500 130.0000 ;
      RECT 227.0500 129.3800 230.7500 130.0000 ;
      RECT 223.0500 129.3800 226.7500 130.0000 ;
      RECT 219.0500 129.3800 222.7500 130.0000 ;
      RECT 215.0500 129.3800 218.7500 130.0000 ;
      RECT 211.0500 129.3800 214.7500 130.0000 ;
      RECT 207.0500 129.3800 210.7500 130.0000 ;
      RECT 203.0500 129.3800 206.7500 130.0000 ;
      RECT 199.0500 129.3800 202.7500 130.0000 ;
      RECT 195.0500 129.3800 198.7500 130.0000 ;
      RECT 191.0500 129.3800 194.7500 130.0000 ;
      RECT 187.0500 129.3800 190.7500 130.0000 ;
      RECT 183.0500 129.3800 186.7500 130.0000 ;
      RECT 179.0500 129.3800 182.7500 130.0000 ;
      RECT 175.0500 129.3800 178.7500 130.0000 ;
      RECT 171.0500 129.3800 174.7500 130.0000 ;
      RECT 167.0500 129.3800 170.7500 130.0000 ;
      RECT 163.0500 129.3800 166.7500 130.0000 ;
      RECT 159.0500 129.3800 162.7500 130.0000 ;
      RECT 155.0500 129.3800 158.7500 130.0000 ;
      RECT 151.0500 129.3800 154.7500 130.0000 ;
      RECT 147.0500 129.3800 150.7500 130.0000 ;
      RECT 143.0500 129.3800 146.7500 130.0000 ;
      RECT 139.0500 129.3800 142.7500 130.0000 ;
      RECT 135.0500 129.3800 138.7500 130.0000 ;
      RECT 131.0500 129.3800 134.7500 130.0000 ;
      RECT 127.0500 129.3800 130.7500 130.0000 ;
      RECT 123.0500 129.3800 126.7500 130.0000 ;
      RECT 119.0500 129.3800 122.7500 130.0000 ;
      RECT 115.0500 129.3800 118.7500 130.0000 ;
      RECT 111.0500 129.3800 114.7500 130.0000 ;
      RECT 107.0500 129.3800 110.7500 130.0000 ;
      RECT 103.0500 129.3800 106.7500 130.0000 ;
      RECT 99.0500 129.3800 102.7500 130.0000 ;
      RECT 95.0500 129.3800 98.7500 130.0000 ;
      RECT 91.0500 129.3800 94.7500 130.0000 ;
      RECT 87.0500 129.3800 90.7500 130.0000 ;
      RECT 83.0500 129.3800 86.7500 130.0000 ;
      RECT 79.0500 129.3800 82.7500 130.0000 ;
      RECT 75.0500 129.3800 78.7500 130.0000 ;
      RECT 71.0500 129.3800 74.7500 130.0000 ;
      RECT 67.0500 129.3800 70.7500 130.0000 ;
      RECT 63.0500 129.3800 66.7500 130.0000 ;
      RECT 59.0500 129.3800 62.7500 130.0000 ;
      RECT 55.0500 129.3800 58.7500 130.0000 ;
      RECT 51.0500 129.3800 54.7500 130.0000 ;
      RECT 47.0500 129.3800 50.7500 130.0000 ;
      RECT 0.0000 129.3800 46.7500 130.0000 ;
      RECT 0.0000 115.1600 730.0000 129.3800 ;
      RECT 698.1300 14.8400 698.8100 115.1600 ;
      RECT 682.9000 14.8400 696.8100 115.1600 ;
      RECT 680.9000 14.8400 681.5800 115.1600 ;
      RECT 665.6700 14.8400 679.5800 115.1600 ;
      RECT 663.6700 14.8400 664.3500 115.1600 ;
      RECT 648.4400 14.8400 662.3500 115.1600 ;
      RECT 646.4400 14.8400 647.1200 115.1600 ;
      RECT 631.2100 14.8400 645.1200 115.1600 ;
      RECT 629.2100 14.8400 629.8900 115.1600 ;
      RECT 613.9800 14.8400 627.8900 115.1600 ;
      RECT 611.9800 14.8400 612.6600 115.1600 ;
      RECT 596.7500 14.8400 610.6600 115.1600 ;
      RECT 594.7500 14.8400 595.4300 115.1600 ;
      RECT 579.5200 14.8400 593.4300 115.1600 ;
      RECT 577.5200 14.8400 578.2000 115.1600 ;
      RECT 562.2900 14.8400 576.2000 115.1600 ;
      RECT 560.2900 14.8400 560.9700 115.1600 ;
      RECT 545.0600 14.8400 558.9700 115.1600 ;
      RECT 543.0600 14.8400 543.7400 115.1600 ;
      RECT 527.8300 14.8400 541.7400 115.1600 ;
      RECT 525.8300 14.8400 526.5100 115.1600 ;
      RECT 510.6000 14.8400 524.5100 115.1600 ;
      RECT 508.6000 14.8400 509.2800 115.1600 ;
      RECT 493.3700 14.8400 507.2800 115.1600 ;
      RECT 491.3700 14.8400 492.0500 115.1600 ;
      RECT 476.1400 14.8400 490.0500 115.1600 ;
      RECT 474.1400 14.8400 474.8200 115.1600 ;
      RECT 458.9100 14.8400 472.8200 115.1600 ;
      RECT 456.9100 14.8400 457.5900 115.1600 ;
      RECT 441.6800 14.8400 455.5900 115.1600 ;
      RECT 439.6800 14.8400 440.3600 115.1600 ;
      RECT 424.4500 14.8400 438.3600 115.1600 ;
      RECT 422.4500 14.8400 423.1300 115.1600 ;
      RECT 407.2200 14.8400 421.1300 115.1600 ;
      RECT 405.2200 14.8400 405.9000 115.1600 ;
      RECT 389.9900 14.8400 403.9000 115.1600 ;
      RECT 387.9900 14.8400 388.6700 115.1600 ;
      RECT 372.7600 14.8400 386.6700 115.1600 ;
      RECT 370.7600 14.8400 371.4400 115.1600 ;
      RECT 355.5300 14.8400 369.4400 115.1600 ;
      RECT 353.5300 14.8400 354.2100 115.1600 ;
      RECT 338.3000 14.8400 352.2100 115.1600 ;
      RECT 336.3000 14.8400 336.9800 115.1600 ;
      RECT 321.0700 14.8400 334.9800 115.1600 ;
      RECT 319.0700 14.8400 319.7500 115.1600 ;
      RECT 303.8400 14.8400 317.7500 115.1600 ;
      RECT 301.8400 14.8400 302.5200 115.1600 ;
      RECT 286.6100 14.8400 300.5200 115.1600 ;
      RECT 284.6100 14.8400 285.2900 115.1600 ;
      RECT 269.3800 14.8400 283.2900 115.1600 ;
      RECT 267.3800 14.8400 268.0600 115.1600 ;
      RECT 252.1500 14.8400 266.0600 115.1600 ;
      RECT 250.1500 14.8400 250.8300 115.1600 ;
      RECT 234.9200 14.8400 248.8300 115.1600 ;
      RECT 232.9200 14.8400 233.6000 115.1600 ;
      RECT 217.6900 14.8400 231.6000 115.1600 ;
      RECT 215.6900 14.8400 216.3700 115.1600 ;
      RECT 200.4600 14.8400 214.3700 115.1600 ;
      RECT 198.4600 14.8400 199.1400 115.1600 ;
      RECT 183.2300 14.8400 197.1400 115.1600 ;
      RECT 181.2300 14.8400 181.9100 115.1600 ;
      RECT 166.0000 14.8400 179.9100 115.1600 ;
      RECT 164.0000 14.8400 164.6800 115.1600 ;
      RECT 148.7700 14.8400 162.6800 115.1600 ;
      RECT 146.7700 14.8400 147.4500 115.1600 ;
      RECT 131.5400 14.8400 145.4500 115.1600 ;
      RECT 129.5400 14.8400 130.2200 115.1600 ;
      RECT 114.3100 14.8400 128.2200 115.1600 ;
      RECT 112.3100 14.8400 112.9900 115.1600 ;
      RECT 97.0800 14.8400 110.9900 115.1600 ;
      RECT 95.0800 14.8400 95.7600 115.1600 ;
      RECT 79.8500 14.8400 93.7600 115.1600 ;
      RECT 77.8500 14.8400 78.5300 115.1600 ;
      RECT 62.6200 14.8400 76.5300 115.1600 ;
      RECT 60.6200 14.8400 61.3000 115.1600 ;
      RECT 45.3900 14.8400 59.3000 115.1600 ;
      RECT 43.3900 14.8400 44.0700 115.1600 ;
      RECT 28.1600 14.8400 42.0700 115.1600 ;
      RECT 26.1600 14.8400 26.8400 115.1600 ;
      RECT 0.0000 14.8400 24.8400 115.1600 ;
      RECT 700.1300 14.6750 730.0000 115.1600 ;
      RECT 682.9000 14.6750 698.8100 14.8400 ;
      RECT 665.6700 14.6750 681.5800 14.8400 ;
      RECT 648.4400 14.6750 664.3500 14.8400 ;
      RECT 631.2100 14.6750 647.1200 14.8400 ;
      RECT 613.9800 14.6750 629.8900 14.8400 ;
      RECT 596.7500 14.6750 612.6600 14.8400 ;
      RECT 579.5200 14.6750 595.4300 14.8400 ;
      RECT 562.2900 14.6750 578.2000 14.8400 ;
      RECT 545.0600 14.6750 560.9700 14.8400 ;
      RECT 527.8300 14.6750 543.7400 14.8400 ;
      RECT 510.6000 14.6750 526.5100 14.8400 ;
      RECT 493.3700 14.6750 509.2800 14.8400 ;
      RECT 476.1400 14.6750 492.0500 14.8400 ;
      RECT 458.9100 14.6750 474.8200 14.8400 ;
      RECT 441.6800 14.6750 457.5900 14.8400 ;
      RECT 424.4500 14.6750 440.3600 14.8400 ;
      RECT 407.2200 14.6750 423.1300 14.8400 ;
      RECT 389.9900 14.6750 405.9000 14.8400 ;
      RECT 372.7600 14.6750 388.6700 14.8400 ;
      RECT 355.5300 14.6750 371.4400 14.8400 ;
      RECT 338.3000 14.6750 354.2100 14.8400 ;
      RECT 321.0700 14.6750 336.9800 14.8400 ;
      RECT 303.8400 14.6750 319.7500 14.8400 ;
      RECT 286.6100 14.6750 302.5200 14.8400 ;
      RECT 269.3800 14.6750 285.2900 14.8400 ;
      RECT 252.1500 14.6750 268.0600 14.8400 ;
      RECT 234.9200 14.6750 250.8300 14.8400 ;
      RECT 217.6900 14.6750 233.6000 14.8400 ;
      RECT 200.4600 14.6750 216.3700 14.8400 ;
      RECT 183.2300 14.6750 199.1400 14.8400 ;
      RECT 166.0000 14.6750 181.9100 14.8400 ;
      RECT 148.7700 14.6750 164.6800 14.8400 ;
      RECT 131.5400 14.6750 147.4500 14.8400 ;
      RECT 114.3100 14.6750 130.2200 14.8400 ;
      RECT 97.0800 14.6750 112.9900 14.8400 ;
      RECT 79.8500 14.6750 95.7600 14.8400 ;
      RECT 62.6200 14.6750 78.5300 14.8400 ;
      RECT 45.3900 14.6750 61.3000 14.8400 ;
      RECT 28.1600 14.6750 44.0700 14.8400 ;
      RECT 0.0000 14.6750 26.8400 14.8400 ;
      RECT 0.0000 0.6200 730.0000 14.6750 ;
      RECT 683.0500 0.0000 730.0000 0.6200 ;
      RECT 679.0500 0.0000 682.7500 0.6200 ;
      RECT 675.0500 0.0000 678.7500 0.6200 ;
      RECT 671.0500 0.0000 674.7500 0.6200 ;
      RECT 667.0500 0.0000 670.7500 0.6200 ;
      RECT 663.0500 0.0000 666.7500 0.6200 ;
      RECT 659.0500 0.0000 662.7500 0.6200 ;
      RECT 655.0500 0.0000 658.7500 0.6200 ;
      RECT 651.0500 0.0000 654.7500 0.6200 ;
      RECT 647.0500 0.0000 650.7500 0.6200 ;
      RECT 643.0500 0.0000 646.7500 0.6200 ;
      RECT 639.0500 0.0000 642.7500 0.6200 ;
      RECT 635.0500 0.0000 638.7500 0.6200 ;
      RECT 631.0500 0.0000 634.7500 0.6200 ;
      RECT 627.0500 0.0000 630.7500 0.6200 ;
      RECT 623.0500 0.0000 626.7500 0.6200 ;
      RECT 619.0500 0.0000 622.7500 0.6200 ;
      RECT 615.0500 0.0000 618.7500 0.6200 ;
      RECT 611.0500 0.0000 614.7500 0.6200 ;
      RECT 607.0500 0.0000 610.7500 0.6200 ;
      RECT 603.0500 0.0000 606.7500 0.6200 ;
      RECT 599.0500 0.0000 602.7500 0.6200 ;
      RECT 595.0500 0.0000 598.7500 0.6200 ;
      RECT 591.0500 0.0000 594.7500 0.6200 ;
      RECT 587.0500 0.0000 590.7500 0.6200 ;
      RECT 583.0500 0.0000 586.7500 0.6200 ;
      RECT 579.0500 0.0000 582.7500 0.6200 ;
      RECT 575.0500 0.0000 578.7500 0.6200 ;
      RECT 571.0500 0.0000 574.7500 0.6200 ;
      RECT 567.0500 0.0000 570.7500 0.6200 ;
      RECT 563.0500 0.0000 566.7500 0.6200 ;
      RECT 559.0500 0.0000 562.7500 0.6200 ;
      RECT 555.0500 0.0000 558.7500 0.6200 ;
      RECT 551.0500 0.0000 554.7500 0.6200 ;
      RECT 547.0500 0.0000 550.7500 0.6200 ;
      RECT 543.0500 0.0000 546.7500 0.6200 ;
      RECT 539.0500 0.0000 542.7500 0.6200 ;
      RECT 535.0500 0.0000 538.7500 0.6200 ;
      RECT 531.0500 0.0000 534.7500 0.6200 ;
      RECT 527.0500 0.0000 530.7500 0.6200 ;
      RECT 523.0500 0.0000 526.7500 0.6200 ;
      RECT 519.0500 0.0000 522.7500 0.6200 ;
      RECT 515.0500 0.0000 518.7500 0.6200 ;
      RECT 511.0500 0.0000 514.7500 0.6200 ;
      RECT 507.0500 0.0000 510.7500 0.6200 ;
      RECT 503.0500 0.0000 506.7500 0.6200 ;
      RECT 499.0500 0.0000 502.7500 0.6200 ;
      RECT 495.0500 0.0000 498.7500 0.6200 ;
      RECT 491.0500 0.0000 494.7500 0.6200 ;
      RECT 487.0500 0.0000 490.7500 0.6200 ;
      RECT 483.0500 0.0000 486.7500 0.6200 ;
      RECT 479.0500 0.0000 482.7500 0.6200 ;
      RECT 475.0500 0.0000 478.7500 0.6200 ;
      RECT 471.0500 0.0000 474.7500 0.6200 ;
      RECT 467.0500 0.0000 470.7500 0.6200 ;
      RECT 463.0500 0.0000 466.7500 0.6200 ;
      RECT 459.0500 0.0000 462.7500 0.6200 ;
      RECT 455.0500 0.0000 458.7500 0.6200 ;
      RECT 451.0500 0.0000 454.7500 0.6200 ;
      RECT 447.0500 0.0000 450.7500 0.6200 ;
      RECT 443.0500 0.0000 446.7500 0.6200 ;
      RECT 439.0500 0.0000 442.7500 0.6200 ;
      RECT 435.0500 0.0000 438.7500 0.6200 ;
      RECT 431.0500 0.0000 434.7500 0.6200 ;
      RECT 427.0500 0.0000 430.7500 0.6200 ;
      RECT 423.0500 0.0000 426.7500 0.6200 ;
      RECT 419.0500 0.0000 422.7500 0.6200 ;
      RECT 415.0500 0.0000 418.7500 0.6200 ;
      RECT 411.0500 0.0000 414.7500 0.6200 ;
      RECT 407.0500 0.0000 410.7500 0.6200 ;
      RECT 403.0500 0.0000 406.7500 0.6200 ;
      RECT 399.0500 0.0000 402.7500 0.6200 ;
      RECT 395.0500 0.0000 398.7500 0.6200 ;
      RECT 391.0500 0.0000 394.7500 0.6200 ;
      RECT 387.0500 0.0000 390.7500 0.6200 ;
      RECT 383.0500 0.0000 386.7500 0.6200 ;
      RECT 379.0500 0.0000 382.7500 0.6200 ;
      RECT 375.0500 0.0000 378.7500 0.6200 ;
      RECT 371.0500 0.0000 374.7500 0.6200 ;
      RECT 367.0500 0.0000 370.7500 0.6200 ;
      RECT 363.0500 0.0000 366.7500 0.6200 ;
      RECT 359.0500 0.0000 362.7500 0.6200 ;
      RECT 355.0500 0.0000 358.7500 0.6200 ;
      RECT 351.0500 0.0000 354.7500 0.6200 ;
      RECT 347.0500 0.0000 350.7500 0.6200 ;
      RECT 343.0500 0.0000 346.7500 0.6200 ;
      RECT 339.0500 0.0000 342.7500 0.6200 ;
      RECT 335.0500 0.0000 338.7500 0.6200 ;
      RECT 331.0500 0.0000 334.7500 0.6200 ;
      RECT 327.0500 0.0000 330.7500 0.6200 ;
      RECT 323.0500 0.0000 326.7500 0.6200 ;
      RECT 319.0500 0.0000 322.7500 0.6200 ;
      RECT 315.0500 0.0000 318.7500 0.6200 ;
      RECT 311.0500 0.0000 314.7500 0.6200 ;
      RECT 307.0500 0.0000 310.7500 0.6200 ;
      RECT 303.0500 0.0000 306.7500 0.6200 ;
      RECT 299.0500 0.0000 302.7500 0.6200 ;
      RECT 295.0500 0.0000 298.7500 0.6200 ;
      RECT 291.0500 0.0000 294.7500 0.6200 ;
      RECT 287.0500 0.0000 290.7500 0.6200 ;
      RECT 283.0500 0.0000 286.7500 0.6200 ;
      RECT 279.0500 0.0000 282.7500 0.6200 ;
      RECT 275.0500 0.0000 278.7500 0.6200 ;
      RECT 271.0500 0.0000 274.7500 0.6200 ;
      RECT 267.0500 0.0000 270.7500 0.6200 ;
      RECT 263.0500 0.0000 266.7500 0.6200 ;
      RECT 259.0500 0.0000 262.7500 0.6200 ;
      RECT 255.0500 0.0000 258.7500 0.6200 ;
      RECT 251.0500 0.0000 254.7500 0.6200 ;
      RECT 247.0500 0.0000 250.7500 0.6200 ;
      RECT 243.0500 0.0000 246.7500 0.6200 ;
      RECT 239.0500 0.0000 242.7500 0.6200 ;
      RECT 235.0500 0.0000 238.7500 0.6200 ;
      RECT 231.0500 0.0000 234.7500 0.6200 ;
      RECT 227.0500 0.0000 230.7500 0.6200 ;
      RECT 223.0500 0.0000 226.7500 0.6200 ;
      RECT 219.0500 0.0000 222.7500 0.6200 ;
      RECT 215.0500 0.0000 218.7500 0.6200 ;
      RECT 211.0500 0.0000 214.7500 0.6200 ;
      RECT 207.0500 0.0000 210.7500 0.6200 ;
      RECT 203.0500 0.0000 206.7500 0.6200 ;
      RECT 199.0500 0.0000 202.7500 0.6200 ;
      RECT 195.0500 0.0000 198.7500 0.6200 ;
      RECT 191.0500 0.0000 194.7500 0.6200 ;
      RECT 187.0500 0.0000 190.7500 0.6200 ;
      RECT 183.0500 0.0000 186.7500 0.6200 ;
      RECT 179.0500 0.0000 182.7500 0.6200 ;
      RECT 175.0500 0.0000 178.7500 0.6200 ;
      RECT 171.0500 0.0000 174.7500 0.6200 ;
      RECT 167.0500 0.0000 170.7500 0.6200 ;
      RECT 163.0500 0.0000 166.7500 0.6200 ;
      RECT 159.0500 0.0000 162.7500 0.6200 ;
      RECT 155.0500 0.0000 158.7500 0.6200 ;
      RECT 151.0500 0.0000 154.7500 0.6200 ;
      RECT 147.0500 0.0000 150.7500 0.6200 ;
      RECT 143.0500 0.0000 146.7500 0.6200 ;
      RECT 139.0500 0.0000 142.7500 0.6200 ;
      RECT 135.0500 0.0000 138.7500 0.6200 ;
      RECT 131.0500 0.0000 134.7500 0.6200 ;
      RECT 127.0500 0.0000 130.7500 0.6200 ;
      RECT 123.0500 0.0000 126.7500 0.6200 ;
      RECT 119.0500 0.0000 122.7500 0.6200 ;
      RECT 115.0500 0.0000 118.7500 0.6200 ;
      RECT 111.0500 0.0000 114.7500 0.6200 ;
      RECT 107.0500 0.0000 110.7500 0.6200 ;
      RECT 103.0500 0.0000 106.7500 0.6200 ;
      RECT 99.0500 0.0000 102.7500 0.6200 ;
      RECT 95.0500 0.0000 98.7500 0.6200 ;
      RECT 91.0500 0.0000 94.7500 0.6200 ;
      RECT 87.0500 0.0000 90.7500 0.6200 ;
      RECT 83.0500 0.0000 86.7500 0.6200 ;
      RECT 79.0500 0.0000 82.7500 0.6200 ;
      RECT 75.0500 0.0000 78.7500 0.6200 ;
      RECT 71.0500 0.0000 74.7500 0.6200 ;
      RECT 67.0500 0.0000 70.7500 0.6200 ;
      RECT 63.0500 0.0000 66.7500 0.6200 ;
      RECT 59.0500 0.0000 62.7500 0.6200 ;
      RECT 55.0500 0.0000 58.7500 0.6200 ;
      RECT 51.0500 0.0000 54.7500 0.6200 ;
      RECT 47.0500 0.0000 50.7500 0.6200 ;
      RECT 0.0000 0.0000 46.7500 0.6200 ;
  END
END sram_w16_out

END LIBRARY
