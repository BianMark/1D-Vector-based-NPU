##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Thu Mar 20 14:19:58 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16_in
  CLASS BLOCK ;
  SIZE 320.0000 BY 120.0000 ;
  FOREIGN sram_w16_in 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 52.1500 0.5200 52.2500 ;
    END
  END CLK
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 33.8500 0.0000 33.9500 0.5200 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.8500 0.0000 37.9500 0.5200 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 41.8500 0.0000 41.9500 0.5200 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 45.8500 0.0000 45.9500 0.5200 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 49.8500 0.0000 49.9500 0.5200 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 53.8500 0.0000 53.9500 0.5200 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 57.8500 0.0000 57.9500 0.5200 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 61.8500 0.0000 61.9500 0.5200 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 65.8500 0.0000 65.9500 0.5200 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 69.8500 0.0000 69.9500 0.5200 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 73.8500 0.0000 73.9500 0.5200 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 77.8500 0.0000 77.9500 0.5200 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 81.8500 0.0000 81.9500 0.5200 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 85.8500 0.0000 85.9500 0.5200 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 89.8500 0.0000 89.9500 0.5200 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 93.8500 0.0000 93.9500 0.5200 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 97.8500 0.0000 97.9500 0.5200 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 101.8500 0.0000 101.9500 0.5200 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 105.8500 0.0000 105.9500 0.5200 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 109.8500 0.0000 109.9500 0.5200 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 113.8500 0.0000 113.9500 0.5200 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 117.8500 0.0000 117.9500 0.5200 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 121.8500 0.0000 121.9500 0.5200 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 125.8500 0.0000 125.9500 0.5200 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 129.8500 0.0000 129.9500 0.5200 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 133.8500 0.0000 133.9500 0.5200 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 137.8500 0.0000 137.9500 0.5200 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 141.8500 0.0000 141.9500 0.5200 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 145.8500 0.0000 145.9500 0.5200 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 149.8500 0.0000 149.9500 0.5200 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 153.8500 0.0000 153.9500 0.5200 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 157.8500 0.0000 157.9500 0.5200 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 161.8500 0.0000 161.9500 0.5200 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 165.8500 0.0000 165.9500 0.5200 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 169.8500 0.0000 169.9500 0.5200 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 173.8500 0.0000 173.9500 0.5200 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 177.8500 0.0000 177.9500 0.5200 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 181.8500 0.0000 181.9500 0.5200 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 185.8500 0.0000 185.9500 0.5200 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 189.8500 0.0000 189.9500 0.5200 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 193.8500 0.0000 193.9500 0.5200 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 197.8500 0.0000 197.9500 0.5200 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 201.8500 0.0000 201.9500 0.5200 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 205.8500 0.0000 205.9500 0.5200 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 209.8500 0.0000 209.9500 0.5200 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 213.8500 0.0000 213.9500 0.5200 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 217.8500 0.0000 217.9500 0.5200 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 221.8500 0.0000 221.9500 0.5200 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 225.8500 0.0000 225.9500 0.5200 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 229.8500 0.0000 229.9500 0.5200 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 233.8500 0.0000 233.9500 0.5200 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 237.8500 0.0000 237.9500 0.5200 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 241.8500 0.0000 241.9500 0.5200 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 245.8500 0.0000 245.9500 0.5200 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 249.8500 0.0000 249.9500 0.5200 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 253.8500 0.0000 253.9500 0.5200 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 257.8500 0.0000 257.9500 0.5200 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 261.8500 0.0000 261.9500 0.5200 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 265.8500 0.0000 265.9500 0.5200 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 269.8500 0.0000 269.9500 0.5200 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 273.8500 0.0000 273.9500 0.5200 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 277.8500 0.0000 277.9500 0.5200 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 281.8500 0.0000 281.9500 0.5200 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 285.8500 0.0000 285.9500 0.5200 ;
    END
  END D[0]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 33.8500 119.4800 33.9500 120.0000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 37.8500 119.4800 37.9500 120.0000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 41.8500 119.4800 41.9500 120.0000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 45.8500 119.4800 45.9500 120.0000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 49.8500 119.4800 49.9500 120.0000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 53.8500 119.4800 53.9500 120.0000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 57.8500 119.4800 57.9500 120.0000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 61.8500 119.4800 61.9500 120.0000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 65.8500 119.4800 65.9500 120.0000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 69.8500 119.4800 69.9500 120.0000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 73.8500 119.4800 73.9500 120.0000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 77.8500 119.4800 77.9500 120.0000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 81.8500 119.4800 81.9500 120.0000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 85.8500 119.4800 85.9500 120.0000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 89.8500 119.4800 89.9500 120.0000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 93.8500 119.4800 93.9500 120.0000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 97.8500 119.4800 97.9500 120.0000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 101.8500 119.4800 101.9500 120.0000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 105.8500 119.4800 105.9500 120.0000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 109.8500 119.4800 109.9500 120.0000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 113.8500 119.4800 113.9500 120.0000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 117.8500 119.4800 117.9500 120.0000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 121.8500 119.4800 121.9500 120.0000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 125.8500 119.4800 125.9500 120.0000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 129.8500 119.4800 129.9500 120.0000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 133.8500 119.4800 133.9500 120.0000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 137.8500 119.4800 137.9500 120.0000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 141.8500 119.4800 141.9500 120.0000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 145.8500 119.4800 145.9500 120.0000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 149.8500 119.4800 149.9500 120.0000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 153.8500 119.4800 153.9500 120.0000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 157.8500 119.4800 157.9500 120.0000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 161.8500 119.4800 161.9500 120.0000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 165.8500 119.4800 165.9500 120.0000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 169.8500 119.4800 169.9500 120.0000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 173.8500 119.4800 173.9500 120.0000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 177.8500 119.4800 177.9500 120.0000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 181.8500 119.4800 181.9500 120.0000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 185.8500 119.4800 185.9500 120.0000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 189.8500 119.4800 189.9500 120.0000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 193.8500 119.4800 193.9500 120.0000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 197.8500 119.4800 197.9500 120.0000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 201.8500 119.4800 201.9500 120.0000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 205.8500 119.4800 205.9500 120.0000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 209.8500 119.4800 209.9500 120.0000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 213.8500 119.4800 213.9500 120.0000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 217.8500 119.4800 217.9500 120.0000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 221.8500 119.4800 221.9500 120.0000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 225.8500 119.4800 225.9500 120.0000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 229.8500 119.4800 229.9500 120.0000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 233.8500 119.4800 233.9500 120.0000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 237.8500 119.4800 237.9500 120.0000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 241.8500 119.4800 241.9500 120.0000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 245.8500 119.4800 245.9500 120.0000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 249.8500 119.4800 249.9500 120.0000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 253.8500 119.4800 253.9500 120.0000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 257.8500 119.4800 257.9500 120.0000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 261.8500 119.4800 261.9500 120.0000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 265.8500 119.4800 265.9500 120.0000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 269.8500 119.4800 269.9500 120.0000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 273.8500 119.4800 273.9500 120.0000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 277.8500 119.4800 277.9500 120.0000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 281.8500 119.4800 281.9500 120.0000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 285.8500 119.4800 285.9500 120.0000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 56.1500 0.5200 56.2500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 48.1500 0.5200 48.2500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 72.1500 0.5200 72.2500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 68.1500 0.5200 68.2500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 64.1500 0.5200 64.2500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 60.1500 0.5200 60.2500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 151.1750 10.0000 152.1750 110.0000 ;
        RECT 136.6000 10.0000 137.6000 110.0000 ;
        RECT 122.0250 10.0000 123.0250 110.0000 ;
        RECT 107.4500 10.0000 108.4500 110.0000 ;
        RECT 92.8750 10.0000 93.8750 110.0000 ;
        RECT 78.3000 10.0000 79.3000 110.0000 ;
        RECT 63.7250 10.0000 64.7250 110.0000 ;
        RECT 49.1500 10.0000 50.1500 110.0000 ;
        RECT 34.5750 10.0000 35.5750 110.0000 ;
        RECT 20.0000 10.0000 21.0000 110.0000 ;
        RECT 296.9250 10.0000 297.9250 110.0000 ;
        RECT 282.3500 10.0000 283.3500 110.0000 ;
        RECT 267.7750 10.0000 268.7750 110.0000 ;
        RECT 253.2000 10.0000 254.2000 110.0000 ;
        RECT 238.6250 10.0000 239.6250 110.0000 ;
        RECT 224.0500 10.0000 225.0500 110.0000 ;
        RECT 209.4750 10.0000 210.4750 110.0000 ;
        RECT 194.9000 10.0000 195.9000 110.0000 ;
        RECT 180.3250 10.0000 181.3250 110.0000 ;
        RECT 165.7500 10.0000 166.7500 110.0000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 153.1750 10.0000 154.1750 110.0000 ;
        RECT 138.6000 10.0000 139.6000 110.0000 ;
        RECT 124.0250 10.0000 125.0250 110.0000 ;
        RECT 109.4500 10.0000 110.4500 110.0000 ;
        RECT 94.8750 10.0000 95.8750 110.0000 ;
        RECT 80.3000 10.0000 81.3000 110.0000 ;
        RECT 65.7250 10.0000 66.7250 110.0000 ;
        RECT 51.1500 10.0000 52.1500 110.0000 ;
        RECT 36.5750 10.0000 37.5750 110.0000 ;
        RECT 22.0000 10.0000 23.0000 110.0000 ;
        RECT 167.7500 10.0000 168.7500 110.0000 ;
        RECT 182.3250 10.0000 183.3250 110.0000 ;
        RECT 196.9000 10.0000 197.9000 110.0000 ;
        RECT 211.4750 10.0000 212.4750 110.0000 ;
        RECT 226.0500 10.0000 227.0500 110.0000 ;
        RECT 240.6250 10.0000 241.6250 110.0000 ;
        RECT 255.2000 10.0000 256.2000 110.0000 ;
        RECT 269.7750 10.0000 270.7750 110.0000 ;
        RECT 284.3500 10.0000 285.3500 110.0000 ;
        RECT 298.9250 10.0000 299.9250 110.0000 ;
        RECT 36.5750 9.8350 37.5750 10.1650 ;
        RECT 22.0000 9.8350 23.0000 10.1650 ;
        RECT 51.1500 9.8350 52.1500 10.1650 ;
        RECT 65.7250 9.8350 66.7250 10.1650 ;
        RECT 94.8750 9.8350 95.8750 10.1650 ;
        RECT 80.3000 9.8350 81.3000 10.1650 ;
        RECT 109.4500 9.8350 110.4500 10.1650 ;
        RECT 138.6000 9.8350 139.6000 10.1650 ;
        RECT 124.0250 9.8350 125.0250 10.1650 ;
        RECT 153.1750 9.8350 154.1750 10.1650 ;
        RECT 167.7500 9.8350 168.7500 10.1650 ;
        RECT 196.9000 9.8350 197.9000 10.1650 ;
        RECT 182.3250 9.8350 183.3250 10.1650 ;
        RECT 211.4750 9.8350 212.4750 10.1650 ;
        RECT 226.0500 9.8350 227.0500 10.1650 ;
        RECT 255.2000 9.8350 256.2000 10.1650 ;
        RECT 240.6250 9.8350 241.6250 10.1650 ;
        RECT 269.7750 9.8350 270.7750 10.1650 ;
        RECT 298.9250 9.8350 299.9250 10.1650 ;
        RECT 284.3500 9.8350 285.3500 10.1650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 320.0000 120.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 320.0000 120.0000 ;
    LAYER M3 ;
      RECT 0.0000 72.3500 320.0000 120.0000 ;
      RECT 0.6200 72.0500 320.0000 72.3500 ;
      RECT 0.0000 68.3500 320.0000 72.0500 ;
      RECT 0.6200 68.0500 320.0000 68.3500 ;
      RECT 0.0000 64.3500 320.0000 68.0500 ;
      RECT 0.6200 64.0500 320.0000 64.3500 ;
      RECT 0.0000 60.3500 320.0000 64.0500 ;
      RECT 0.6200 60.0500 320.0000 60.3500 ;
      RECT 0.0000 56.3500 320.0000 60.0500 ;
      RECT 0.6200 56.0500 320.0000 56.3500 ;
      RECT 0.0000 52.3500 320.0000 56.0500 ;
      RECT 0.6200 52.0500 320.0000 52.3500 ;
      RECT 0.0000 48.3500 320.0000 52.0500 ;
      RECT 0.6200 48.0500 320.0000 48.3500 ;
      RECT 0.0000 0.0000 320.0000 48.0500 ;
    LAYER M4 ;
      RECT 286.0500 119.3800 320.0000 120.0000 ;
      RECT 282.0500 119.3800 285.7500 120.0000 ;
      RECT 278.0500 119.3800 281.7500 120.0000 ;
      RECT 274.0500 119.3800 277.7500 120.0000 ;
      RECT 270.0500 119.3800 273.7500 120.0000 ;
      RECT 266.0500 119.3800 269.7500 120.0000 ;
      RECT 262.0500 119.3800 265.7500 120.0000 ;
      RECT 258.0500 119.3800 261.7500 120.0000 ;
      RECT 254.0500 119.3800 257.7500 120.0000 ;
      RECT 250.0500 119.3800 253.7500 120.0000 ;
      RECT 246.0500 119.3800 249.7500 120.0000 ;
      RECT 242.0500 119.3800 245.7500 120.0000 ;
      RECT 238.0500 119.3800 241.7500 120.0000 ;
      RECT 234.0500 119.3800 237.7500 120.0000 ;
      RECT 230.0500 119.3800 233.7500 120.0000 ;
      RECT 226.0500 119.3800 229.7500 120.0000 ;
      RECT 222.0500 119.3800 225.7500 120.0000 ;
      RECT 218.0500 119.3800 221.7500 120.0000 ;
      RECT 214.0500 119.3800 217.7500 120.0000 ;
      RECT 210.0500 119.3800 213.7500 120.0000 ;
      RECT 206.0500 119.3800 209.7500 120.0000 ;
      RECT 202.0500 119.3800 205.7500 120.0000 ;
      RECT 198.0500 119.3800 201.7500 120.0000 ;
      RECT 194.0500 119.3800 197.7500 120.0000 ;
      RECT 190.0500 119.3800 193.7500 120.0000 ;
      RECT 186.0500 119.3800 189.7500 120.0000 ;
      RECT 182.0500 119.3800 185.7500 120.0000 ;
      RECT 178.0500 119.3800 181.7500 120.0000 ;
      RECT 174.0500 119.3800 177.7500 120.0000 ;
      RECT 170.0500 119.3800 173.7500 120.0000 ;
      RECT 166.0500 119.3800 169.7500 120.0000 ;
      RECT 162.0500 119.3800 165.7500 120.0000 ;
      RECT 158.0500 119.3800 161.7500 120.0000 ;
      RECT 154.0500 119.3800 157.7500 120.0000 ;
      RECT 150.0500 119.3800 153.7500 120.0000 ;
      RECT 146.0500 119.3800 149.7500 120.0000 ;
      RECT 142.0500 119.3800 145.7500 120.0000 ;
      RECT 138.0500 119.3800 141.7500 120.0000 ;
      RECT 134.0500 119.3800 137.7500 120.0000 ;
      RECT 130.0500 119.3800 133.7500 120.0000 ;
      RECT 126.0500 119.3800 129.7500 120.0000 ;
      RECT 122.0500 119.3800 125.7500 120.0000 ;
      RECT 118.0500 119.3800 121.7500 120.0000 ;
      RECT 114.0500 119.3800 117.7500 120.0000 ;
      RECT 110.0500 119.3800 113.7500 120.0000 ;
      RECT 106.0500 119.3800 109.7500 120.0000 ;
      RECT 102.0500 119.3800 105.7500 120.0000 ;
      RECT 98.0500 119.3800 101.7500 120.0000 ;
      RECT 94.0500 119.3800 97.7500 120.0000 ;
      RECT 90.0500 119.3800 93.7500 120.0000 ;
      RECT 86.0500 119.3800 89.7500 120.0000 ;
      RECT 82.0500 119.3800 85.7500 120.0000 ;
      RECT 78.0500 119.3800 81.7500 120.0000 ;
      RECT 74.0500 119.3800 77.7500 120.0000 ;
      RECT 70.0500 119.3800 73.7500 120.0000 ;
      RECT 66.0500 119.3800 69.7500 120.0000 ;
      RECT 62.0500 119.3800 65.7500 120.0000 ;
      RECT 58.0500 119.3800 61.7500 120.0000 ;
      RECT 54.0500 119.3800 57.7500 120.0000 ;
      RECT 50.0500 119.3800 53.7500 120.0000 ;
      RECT 46.0500 119.3800 49.7500 120.0000 ;
      RECT 42.0500 119.3800 45.7500 120.0000 ;
      RECT 38.0500 119.3800 41.7500 120.0000 ;
      RECT 34.0500 119.3800 37.7500 120.0000 ;
      RECT 0.0000 119.3800 33.7500 120.0000 ;
      RECT 0.0000 110.1600 320.0000 119.3800 ;
      RECT 298.0850 9.8400 298.7650 110.1600 ;
      RECT 285.5100 9.8400 296.7650 110.1600 ;
      RECT 283.5100 9.8400 284.1900 110.1600 ;
      RECT 270.9350 9.8400 282.1900 110.1600 ;
      RECT 268.9350 9.8400 269.6150 110.1600 ;
      RECT 256.3600 9.8400 267.6150 110.1600 ;
      RECT 254.3600 9.8400 255.0400 110.1600 ;
      RECT 241.7850 9.8400 253.0400 110.1600 ;
      RECT 239.7850 9.8400 240.4650 110.1600 ;
      RECT 227.2100 9.8400 238.4650 110.1600 ;
      RECT 225.2100 9.8400 225.8900 110.1600 ;
      RECT 212.6350 9.8400 223.8900 110.1600 ;
      RECT 210.6350 9.8400 211.3150 110.1600 ;
      RECT 198.0600 9.8400 209.3150 110.1600 ;
      RECT 196.0600 9.8400 196.7400 110.1600 ;
      RECT 183.4850 9.8400 194.7400 110.1600 ;
      RECT 181.4850 9.8400 182.1650 110.1600 ;
      RECT 168.9100 9.8400 180.1650 110.1600 ;
      RECT 166.9100 9.8400 167.5900 110.1600 ;
      RECT 154.3350 9.8400 165.5900 110.1600 ;
      RECT 152.3350 9.8400 153.0150 110.1600 ;
      RECT 139.7600 9.8400 151.0150 110.1600 ;
      RECT 137.7600 9.8400 138.4400 110.1600 ;
      RECT 125.1850 9.8400 136.4400 110.1600 ;
      RECT 123.1850 9.8400 123.8650 110.1600 ;
      RECT 110.6100 9.8400 121.8650 110.1600 ;
      RECT 108.6100 9.8400 109.2900 110.1600 ;
      RECT 96.0350 9.8400 107.2900 110.1600 ;
      RECT 94.0350 9.8400 94.7150 110.1600 ;
      RECT 81.4600 9.8400 92.7150 110.1600 ;
      RECT 79.4600 9.8400 80.1400 110.1600 ;
      RECT 66.8850 9.8400 78.1400 110.1600 ;
      RECT 64.8850 9.8400 65.5650 110.1600 ;
      RECT 52.3100 9.8400 63.5650 110.1600 ;
      RECT 50.3100 9.8400 50.9900 110.1600 ;
      RECT 37.7350 9.8400 48.9900 110.1600 ;
      RECT 35.7350 9.8400 36.4150 110.1600 ;
      RECT 23.1600 9.8400 34.4150 110.1600 ;
      RECT 21.1600 9.8400 21.8400 110.1600 ;
      RECT 0.0000 9.8400 19.8400 110.1600 ;
      RECT 300.0850 9.6750 320.0000 110.1600 ;
      RECT 285.5100 9.6750 298.7650 9.8400 ;
      RECT 270.9350 9.6750 284.1900 9.8400 ;
      RECT 256.3600 9.6750 269.6150 9.8400 ;
      RECT 241.7850 9.6750 255.0400 9.8400 ;
      RECT 227.2100 9.6750 240.4650 9.8400 ;
      RECT 212.6350 9.6750 225.8900 9.8400 ;
      RECT 198.0600 9.6750 211.3150 9.8400 ;
      RECT 183.4850 9.6750 196.7400 9.8400 ;
      RECT 168.9100 9.6750 182.1650 9.8400 ;
      RECT 154.3350 9.6750 167.5900 9.8400 ;
      RECT 139.7600 9.6750 153.0150 9.8400 ;
      RECT 125.1850 9.6750 138.4400 9.8400 ;
      RECT 110.6100 9.6750 123.8650 9.8400 ;
      RECT 96.0350 9.6750 109.2900 9.8400 ;
      RECT 81.4600 9.6750 94.7150 9.8400 ;
      RECT 66.8850 9.6750 80.1400 9.8400 ;
      RECT 52.3100 9.6750 65.5650 9.8400 ;
      RECT 37.7350 9.6750 50.9900 9.8400 ;
      RECT 23.1600 9.6750 36.4150 9.8400 ;
      RECT 0.0000 9.6750 21.8400 9.8400 ;
      RECT 0.0000 0.6200 320.0000 9.6750 ;
      RECT 286.0500 0.0000 320.0000 0.6200 ;
      RECT 282.0500 0.0000 285.7500 0.6200 ;
      RECT 278.0500 0.0000 281.7500 0.6200 ;
      RECT 274.0500 0.0000 277.7500 0.6200 ;
      RECT 270.0500 0.0000 273.7500 0.6200 ;
      RECT 266.0500 0.0000 269.7500 0.6200 ;
      RECT 262.0500 0.0000 265.7500 0.6200 ;
      RECT 258.0500 0.0000 261.7500 0.6200 ;
      RECT 254.0500 0.0000 257.7500 0.6200 ;
      RECT 250.0500 0.0000 253.7500 0.6200 ;
      RECT 246.0500 0.0000 249.7500 0.6200 ;
      RECT 242.0500 0.0000 245.7500 0.6200 ;
      RECT 238.0500 0.0000 241.7500 0.6200 ;
      RECT 234.0500 0.0000 237.7500 0.6200 ;
      RECT 230.0500 0.0000 233.7500 0.6200 ;
      RECT 226.0500 0.0000 229.7500 0.6200 ;
      RECT 222.0500 0.0000 225.7500 0.6200 ;
      RECT 218.0500 0.0000 221.7500 0.6200 ;
      RECT 214.0500 0.0000 217.7500 0.6200 ;
      RECT 210.0500 0.0000 213.7500 0.6200 ;
      RECT 206.0500 0.0000 209.7500 0.6200 ;
      RECT 202.0500 0.0000 205.7500 0.6200 ;
      RECT 198.0500 0.0000 201.7500 0.6200 ;
      RECT 194.0500 0.0000 197.7500 0.6200 ;
      RECT 190.0500 0.0000 193.7500 0.6200 ;
      RECT 186.0500 0.0000 189.7500 0.6200 ;
      RECT 182.0500 0.0000 185.7500 0.6200 ;
      RECT 178.0500 0.0000 181.7500 0.6200 ;
      RECT 174.0500 0.0000 177.7500 0.6200 ;
      RECT 170.0500 0.0000 173.7500 0.6200 ;
      RECT 166.0500 0.0000 169.7500 0.6200 ;
      RECT 162.0500 0.0000 165.7500 0.6200 ;
      RECT 158.0500 0.0000 161.7500 0.6200 ;
      RECT 154.0500 0.0000 157.7500 0.6200 ;
      RECT 150.0500 0.0000 153.7500 0.6200 ;
      RECT 146.0500 0.0000 149.7500 0.6200 ;
      RECT 142.0500 0.0000 145.7500 0.6200 ;
      RECT 138.0500 0.0000 141.7500 0.6200 ;
      RECT 134.0500 0.0000 137.7500 0.6200 ;
      RECT 130.0500 0.0000 133.7500 0.6200 ;
      RECT 126.0500 0.0000 129.7500 0.6200 ;
      RECT 122.0500 0.0000 125.7500 0.6200 ;
      RECT 118.0500 0.0000 121.7500 0.6200 ;
      RECT 114.0500 0.0000 117.7500 0.6200 ;
      RECT 110.0500 0.0000 113.7500 0.6200 ;
      RECT 106.0500 0.0000 109.7500 0.6200 ;
      RECT 102.0500 0.0000 105.7500 0.6200 ;
      RECT 98.0500 0.0000 101.7500 0.6200 ;
      RECT 94.0500 0.0000 97.7500 0.6200 ;
      RECT 90.0500 0.0000 93.7500 0.6200 ;
      RECT 86.0500 0.0000 89.7500 0.6200 ;
      RECT 82.0500 0.0000 85.7500 0.6200 ;
      RECT 78.0500 0.0000 81.7500 0.6200 ;
      RECT 74.0500 0.0000 77.7500 0.6200 ;
      RECT 70.0500 0.0000 73.7500 0.6200 ;
      RECT 66.0500 0.0000 69.7500 0.6200 ;
      RECT 62.0500 0.0000 65.7500 0.6200 ;
      RECT 58.0500 0.0000 61.7500 0.6200 ;
      RECT 54.0500 0.0000 57.7500 0.6200 ;
      RECT 50.0500 0.0000 53.7500 0.6200 ;
      RECT 46.0500 0.0000 49.7500 0.6200 ;
      RECT 42.0500 0.0000 45.7500 0.6200 ;
      RECT 38.0500 0.0000 41.7500 0.6200 ;
      RECT 34.0500 0.0000 37.7500 0.6200 ;
      RECT 0.0000 0.0000 33.7500 0.6200 ;
  END
END sram_w16_in

END LIBRARY
