##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Thu Mar 20 11:53:42 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO core
  CLASS BLOCK ;
  SIZE 524.2000 BY 524.0000 ;
  FOREIGN core 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 97.7500 0.5200 97.8500 ;
    END
  END clk
  PIN sum_out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 84.1500 524.2000 84.2500 ;
    END
  END sum_out[23]
  PIN sum_out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 81.5500 524.2000 81.6500 ;
    END
  END sum_out[22]
  PIN sum_out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 78.9500 524.2000 79.0500 ;
    END
  END sum_out[21]
  PIN sum_out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 76.3500 524.2000 76.4500 ;
    END
  END sum_out[20]
  PIN sum_out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 73.7500 524.2000 73.8500 ;
    END
  END sum_out[19]
  PIN sum_out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 71.1500 524.2000 71.2500 ;
    END
  END sum_out[18]
  PIN sum_out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 68.5500 524.2000 68.6500 ;
    END
  END sum_out[17]
  PIN sum_out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 65.9500 524.2000 66.0500 ;
    END
  END sum_out[16]
  PIN sum_out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 63.3500 524.2000 63.4500 ;
    END
  END sum_out[15]
  PIN sum_out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 60.7500 524.2000 60.8500 ;
    END
  END sum_out[14]
  PIN sum_out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 58.1500 524.2000 58.2500 ;
    END
  END sum_out[13]
  PIN sum_out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 55.5500 524.2000 55.6500 ;
    END
  END sum_out[12]
  PIN sum_out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 52.9500 524.2000 53.0500 ;
    END
  END sum_out[11]
  PIN sum_out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 50.3500 524.2000 50.4500 ;
    END
  END sum_out[10]
  PIN sum_out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 47.7500 524.2000 47.8500 ;
    END
  END sum_out[9]
  PIN sum_out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 45.1500 524.2000 45.2500 ;
    END
  END sum_out[8]
  PIN sum_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 42.5500 524.2000 42.6500 ;
    END
  END sum_out[7]
  PIN sum_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 39.9500 524.2000 40.0500 ;
    END
  END sum_out[6]
  PIN sum_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 37.3500 524.2000 37.4500 ;
    END
  END sum_out[5]
  PIN sum_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 34.7500 524.2000 34.8500 ;
    END
  END sum_out[4]
  PIN sum_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 32.1500 524.2000 32.2500 ;
    END
  END sum_out[3]
  PIN sum_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 29.5500 524.2000 29.6500 ;
    END
  END sum_out[2]
  PIN sum_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 26.9500 524.2000 27.0500 ;
    END
  END sum_out[1]
  PIN sum_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 24.3500 524.2000 24.4500 ;
    END
  END sum_out[0]
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 173.7500 0.5200 173.8500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 177.7500 0.5200 177.8500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 181.7500 0.5200 181.8500 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 185.7500 0.5200 185.8500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 189.7500 0.5200 189.8500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 193.7500 0.5200 193.8500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 197.7500 0.5200 197.8500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 201.7500 0.5200 201.8500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 205.7500 0.5200 205.8500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 209.7500 0.5200 209.8500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 213.7500 0.5200 213.8500 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 217.7500 0.5200 217.8500 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 221.7500 0.5200 221.8500 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 225.7500 0.5200 225.8500 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 229.7500 0.5200 229.8500 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 233.7500 0.5200 233.8500 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 237.7500 0.5200 237.8500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 241.7500 0.5200 241.8500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 245.7500 0.5200 245.8500 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 249.7500 0.5200 249.8500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 253.7500 0.5200 253.8500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 257.7500 0.5200 257.8500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 261.7500 0.5200 261.8500 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 265.7500 0.5200 265.8500 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 269.7500 0.5200 269.8500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 273.7500 0.5200 273.8500 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 277.7500 0.5200 277.8500 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 281.7500 0.5200 281.8500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 285.7500 0.5200 285.8500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 289.7500 0.5200 289.8500 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 293.7500 0.5200 293.8500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 297.7500 0.5200 297.8500 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 301.7500 0.5200 301.8500 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 305.7500 0.5200 305.8500 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 309.7500 0.5200 309.8500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 313.7500 0.5200 313.8500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 317.7500 0.5200 317.8500 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 321.7500 0.5200 321.8500 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 325.7500 0.5200 325.8500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 329.7500 0.5200 329.8500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 333.7500 0.5200 333.8500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 337.7500 0.5200 337.8500 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 341.7500 0.5200 341.8500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 345.7500 0.5200 345.8500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 349.7500 0.5200 349.8500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 353.7500 0.5200 353.8500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 357.7500 0.5200 357.8500 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 361.7500 0.5200 361.8500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 365.7500 0.5200 365.8500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 369.7500 0.5200 369.8500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 373.7500 0.5200 373.8500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 377.7500 0.5200 377.8500 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 381.7500 0.5200 381.8500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 385.7500 0.5200 385.8500 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 389.7500 0.5200 389.8500 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 393.7500 0.5200 393.8500 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 397.7500 0.5200 397.8500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 401.7500 0.5200 401.8500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 405.7500 0.5200 405.8500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 409.7500 0.5200 409.8500 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 413.7500 0.5200 413.8500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 417.7500 0.5200 417.8500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 421.7500 0.5200 421.8500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 425.7500 0.5200 425.8500 ;
    END
  END mem_in[0]
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 500.1500 524.2000 500.2500 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 497.5500 524.2000 497.6500 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 494.9500 524.2000 495.0500 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 492.3500 524.2000 492.4500 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 489.7500 524.2000 489.8500 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 487.1500 524.2000 487.2500 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 484.5500 524.2000 484.6500 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 481.9500 524.2000 482.0500 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 479.3500 524.2000 479.4500 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 476.7500 524.2000 476.8500 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 474.1500 524.2000 474.2500 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 471.5500 524.2000 471.6500 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 468.9500 524.2000 469.0500 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 466.3500 524.2000 466.4500 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 463.7500 524.2000 463.8500 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 461.1500 524.2000 461.2500 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 458.5500 524.2000 458.6500 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 455.9500 524.2000 456.0500 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 453.3500 524.2000 453.4500 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 450.7500 524.2000 450.8500 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 448.1500 524.2000 448.2500 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 445.5500 524.2000 445.6500 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 442.9500 524.2000 443.0500 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 440.3500 524.2000 440.4500 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 437.7500 524.2000 437.8500 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 435.1500 524.2000 435.2500 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 432.5500 524.2000 432.6500 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 429.9500 524.2000 430.0500 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 427.3500 524.2000 427.4500 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 424.7500 524.2000 424.8500 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 422.1500 524.2000 422.2500 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 419.5500 524.2000 419.6500 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 416.9500 524.2000 417.0500 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 414.3500 524.2000 414.4500 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 411.7500 524.2000 411.8500 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 409.1500 524.2000 409.2500 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 406.5500 524.2000 406.6500 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 403.9500 524.2000 404.0500 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 401.3500 524.2000 401.4500 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 398.7500 524.2000 398.8500 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 396.1500 524.2000 396.2500 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 393.5500 524.2000 393.6500 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 390.9500 524.2000 391.0500 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 388.3500 524.2000 388.4500 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 385.7500 524.2000 385.8500 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 383.1500 524.2000 383.2500 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 380.5500 524.2000 380.6500 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 377.9500 524.2000 378.0500 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 375.3500 524.2000 375.4500 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 372.7500 524.2000 372.8500 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 370.1500 524.2000 370.2500 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 367.5500 524.2000 367.6500 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 364.9500 524.2000 365.0500 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 362.3500 524.2000 362.4500 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 359.7500 524.2000 359.8500 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 357.1500 524.2000 357.2500 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 354.5500 524.2000 354.6500 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 351.9500 524.2000 352.0500 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 349.3500 524.2000 349.4500 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 346.7500 524.2000 346.8500 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 344.1500 524.2000 344.2500 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 341.5500 524.2000 341.6500 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 338.9500 524.2000 339.0500 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 336.3500 524.2000 336.4500 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 333.7500 524.2000 333.8500 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 331.1500 524.2000 331.2500 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 328.5500 524.2000 328.6500 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 325.9500 524.2000 326.0500 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 323.3500 524.2000 323.4500 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 320.7500 524.2000 320.8500 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 318.1500 524.2000 318.2500 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 315.5500 524.2000 315.6500 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 312.9500 524.2000 313.0500 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 310.3500 524.2000 310.4500 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 307.7500 524.2000 307.8500 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 305.1500 524.2000 305.2500 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 302.5500 524.2000 302.6500 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 299.9500 524.2000 300.0500 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 297.3500 524.2000 297.4500 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 294.7500 524.2000 294.8500 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 292.1500 524.2000 292.2500 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 289.5500 524.2000 289.6500 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 286.9500 524.2000 287.0500 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 284.3500 524.2000 284.4500 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 281.7500 524.2000 281.8500 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 279.1500 524.2000 279.2500 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 276.5500 524.2000 276.6500 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 273.9500 524.2000 274.0500 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 271.3500 524.2000 271.4500 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 268.7500 524.2000 268.8500 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 266.1500 524.2000 266.2500 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 263.5500 524.2000 263.6500 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 260.9500 524.2000 261.0500 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 258.3500 524.2000 258.4500 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 255.7500 524.2000 255.8500 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 253.1500 524.2000 253.2500 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 250.5500 524.2000 250.6500 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 247.9500 524.2000 248.0500 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 245.3500 524.2000 245.4500 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 242.7500 524.2000 242.8500 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 240.1500 524.2000 240.2500 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 237.5500 524.2000 237.6500 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 234.9500 524.2000 235.0500 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 232.3500 524.2000 232.4500 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 229.7500 524.2000 229.8500 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 227.1500 524.2000 227.2500 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 224.5500 524.2000 224.6500 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 221.9500 524.2000 222.0500 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 219.3500 524.2000 219.4500 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 216.7500 524.2000 216.8500 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 214.1500 524.2000 214.2500 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 211.5500 524.2000 211.6500 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 208.9500 524.2000 209.0500 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 206.3500 524.2000 206.4500 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 203.7500 524.2000 203.8500 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 201.1500 524.2000 201.2500 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 198.5500 524.2000 198.6500 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 195.9500 524.2000 196.0500 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 193.3500 524.2000 193.4500 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 190.7500 524.2000 190.8500 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 188.1500 524.2000 188.2500 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 185.5500 524.2000 185.6500 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 182.9500 524.2000 183.0500 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 180.3500 524.2000 180.4500 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 177.7500 524.2000 177.8500 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 175.1500 524.2000 175.2500 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 172.5500 524.2000 172.6500 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 169.9500 524.2000 170.0500 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 167.3500 524.2000 167.4500 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 164.7500 524.2000 164.8500 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 162.1500 524.2000 162.2500 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 159.5500 524.2000 159.6500 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 156.9500 524.2000 157.0500 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 154.3500 524.2000 154.4500 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 151.7500 524.2000 151.8500 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 149.1500 524.2000 149.2500 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 146.5500 524.2000 146.6500 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 143.9500 524.2000 144.0500 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 141.3500 524.2000 141.4500 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 138.7500 524.2000 138.8500 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 136.1500 524.2000 136.2500 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 133.5500 524.2000 133.6500 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 130.9500 524.2000 131.0500 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 128.3500 524.2000 128.4500 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 125.7500 524.2000 125.8500 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 123.1500 524.2000 123.2500 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 120.5500 524.2000 120.6500 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 117.9500 524.2000 118.0500 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 115.3500 524.2000 115.4500 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 112.7500 524.2000 112.8500 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 110.1500 524.2000 110.2500 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 107.5500 524.2000 107.6500 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 104.9500 524.2000 105.0500 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 102.3500 524.2000 102.4500 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 99.7500 524.2000 99.8500 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 97.1500 524.2000 97.2500 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 94.5500 524.2000 94.6500 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 91.9500 524.2000 92.0500 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 89.3500 524.2000 89.4500 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 523.6800 86.7500 524.2000 86.8500 ;
    END
  END out[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 101.7500 0.5200 101.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 105.7500 0.5200 105.8500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 109.7500 0.5200 109.8500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 113.7500 0.5200 113.8500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 117.7500 0.5200 117.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 121.7500 0.5200 121.8500 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 125.7500 0.5200 125.8500 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 129.7500 0.5200 129.8500 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 133.7500 0.5200 133.8500 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 137.7500 0.5200 137.8500 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 141.7500 0.5200 141.8500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 145.7500 0.5200 145.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 149.7500 0.5200 149.8500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 153.7500 0.5200 153.8500 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 157.7500 0.5200 157.8500 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 161.7500 0.5200 161.8500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 165.7500 0.5200 165.8500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 169.7500 0.5200 169.8500 ;
    END
  END reset
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 524.2000 524.0000 ;
    LAYER M2 ;
      RECT 0.0000 0.0000 524.2000 524.0000 ;
    LAYER M3 ;
      RECT 0.0000 500.3500 524.2000 524.0000 ;
      RECT 0.0000 500.0500 523.5800 500.3500 ;
      RECT 0.0000 497.7500 524.2000 500.0500 ;
      RECT 0.0000 497.4500 523.5800 497.7500 ;
      RECT 0.0000 495.1500 524.2000 497.4500 ;
      RECT 0.0000 494.8500 523.5800 495.1500 ;
      RECT 0.0000 492.5500 524.2000 494.8500 ;
      RECT 0.0000 492.2500 523.5800 492.5500 ;
      RECT 0.0000 489.9500 524.2000 492.2500 ;
      RECT 0.0000 489.6500 523.5800 489.9500 ;
      RECT 0.0000 487.3500 524.2000 489.6500 ;
      RECT 0.0000 487.0500 523.5800 487.3500 ;
      RECT 0.0000 484.7500 524.2000 487.0500 ;
      RECT 0.0000 484.4500 523.5800 484.7500 ;
      RECT 0.0000 482.1500 524.2000 484.4500 ;
      RECT 0.0000 481.8500 523.5800 482.1500 ;
      RECT 0.0000 479.5500 524.2000 481.8500 ;
      RECT 0.0000 479.2500 523.5800 479.5500 ;
      RECT 0.0000 476.9500 524.2000 479.2500 ;
      RECT 0.0000 476.6500 523.5800 476.9500 ;
      RECT 0.0000 474.3500 524.2000 476.6500 ;
      RECT 0.0000 474.0500 523.5800 474.3500 ;
      RECT 0.0000 471.7500 524.2000 474.0500 ;
      RECT 0.0000 471.4500 523.5800 471.7500 ;
      RECT 0.0000 469.1500 524.2000 471.4500 ;
      RECT 0.0000 468.8500 523.5800 469.1500 ;
      RECT 0.0000 466.5500 524.2000 468.8500 ;
      RECT 0.0000 466.2500 523.5800 466.5500 ;
      RECT 0.0000 463.9500 524.2000 466.2500 ;
      RECT 0.0000 463.6500 523.5800 463.9500 ;
      RECT 0.0000 461.3500 524.2000 463.6500 ;
      RECT 0.0000 461.0500 523.5800 461.3500 ;
      RECT 0.0000 458.7500 524.2000 461.0500 ;
      RECT 0.0000 458.4500 523.5800 458.7500 ;
      RECT 0.0000 456.1500 524.2000 458.4500 ;
      RECT 0.0000 455.8500 523.5800 456.1500 ;
      RECT 0.0000 453.5500 524.2000 455.8500 ;
      RECT 0.0000 453.2500 523.5800 453.5500 ;
      RECT 0.0000 450.9500 524.2000 453.2500 ;
      RECT 0.0000 450.6500 523.5800 450.9500 ;
      RECT 0.0000 448.3500 524.2000 450.6500 ;
      RECT 0.0000 448.0500 523.5800 448.3500 ;
      RECT 0.0000 445.7500 524.2000 448.0500 ;
      RECT 0.0000 445.4500 523.5800 445.7500 ;
      RECT 0.0000 443.1500 524.2000 445.4500 ;
      RECT 0.0000 442.8500 523.5800 443.1500 ;
      RECT 0.0000 440.5500 524.2000 442.8500 ;
      RECT 0.0000 440.2500 523.5800 440.5500 ;
      RECT 0.0000 437.9500 524.2000 440.2500 ;
      RECT 0.0000 437.6500 523.5800 437.9500 ;
      RECT 0.0000 435.3500 524.2000 437.6500 ;
      RECT 0.0000 435.0500 523.5800 435.3500 ;
      RECT 0.0000 432.7500 524.2000 435.0500 ;
      RECT 0.0000 432.4500 523.5800 432.7500 ;
      RECT 0.0000 430.1500 524.2000 432.4500 ;
      RECT 0.0000 429.8500 523.5800 430.1500 ;
      RECT 0.0000 427.5500 524.2000 429.8500 ;
      RECT 0.0000 427.2500 523.5800 427.5500 ;
      RECT 0.0000 425.9500 524.2000 427.2500 ;
      RECT 0.6200 425.6500 524.2000 425.9500 ;
      RECT 0.0000 424.9500 524.2000 425.6500 ;
      RECT 0.0000 424.6500 523.5800 424.9500 ;
      RECT 0.0000 422.3500 524.2000 424.6500 ;
      RECT 0.0000 422.0500 523.5800 422.3500 ;
      RECT 0.0000 421.9500 524.2000 422.0500 ;
      RECT 0.6200 421.6500 524.2000 421.9500 ;
      RECT 0.0000 419.7500 524.2000 421.6500 ;
      RECT 0.0000 419.4500 523.5800 419.7500 ;
      RECT 0.0000 417.9500 524.2000 419.4500 ;
      RECT 0.6200 417.6500 524.2000 417.9500 ;
      RECT 0.0000 417.1500 524.2000 417.6500 ;
      RECT 0.0000 416.8500 523.5800 417.1500 ;
      RECT 0.0000 414.5500 524.2000 416.8500 ;
      RECT 0.0000 414.2500 523.5800 414.5500 ;
      RECT 0.0000 413.9500 524.2000 414.2500 ;
      RECT 0.6200 413.6500 524.2000 413.9500 ;
      RECT 0.0000 411.9500 524.2000 413.6500 ;
      RECT 0.0000 411.6500 523.5800 411.9500 ;
      RECT 0.0000 409.9500 524.2000 411.6500 ;
      RECT 0.6200 409.6500 524.2000 409.9500 ;
      RECT 0.0000 409.3500 524.2000 409.6500 ;
      RECT 0.0000 409.0500 523.5800 409.3500 ;
      RECT 0.0000 406.7500 524.2000 409.0500 ;
      RECT 0.0000 406.4500 523.5800 406.7500 ;
      RECT 0.0000 405.9500 524.2000 406.4500 ;
      RECT 0.6200 405.6500 524.2000 405.9500 ;
      RECT 0.0000 404.1500 524.2000 405.6500 ;
      RECT 0.0000 403.8500 523.5800 404.1500 ;
      RECT 0.0000 401.9500 524.2000 403.8500 ;
      RECT 0.6200 401.6500 524.2000 401.9500 ;
      RECT 0.0000 401.5500 524.2000 401.6500 ;
      RECT 0.0000 401.2500 523.5800 401.5500 ;
      RECT 0.0000 398.9500 524.2000 401.2500 ;
      RECT 0.0000 398.6500 523.5800 398.9500 ;
      RECT 0.0000 397.9500 524.2000 398.6500 ;
      RECT 0.6200 397.6500 524.2000 397.9500 ;
      RECT 0.0000 396.3500 524.2000 397.6500 ;
      RECT 0.0000 396.0500 523.5800 396.3500 ;
      RECT 0.0000 393.9500 524.2000 396.0500 ;
      RECT 0.6200 393.7500 524.2000 393.9500 ;
      RECT 0.6200 393.6500 523.5800 393.7500 ;
      RECT 0.0000 393.4500 523.5800 393.6500 ;
      RECT 0.0000 391.1500 524.2000 393.4500 ;
      RECT 0.0000 390.8500 523.5800 391.1500 ;
      RECT 0.0000 389.9500 524.2000 390.8500 ;
      RECT 0.6200 389.6500 524.2000 389.9500 ;
      RECT 0.0000 388.5500 524.2000 389.6500 ;
      RECT 0.0000 388.2500 523.5800 388.5500 ;
      RECT 0.0000 385.9500 524.2000 388.2500 ;
      RECT 0.6200 385.6500 523.5800 385.9500 ;
      RECT 0.0000 383.3500 524.2000 385.6500 ;
      RECT 0.0000 383.0500 523.5800 383.3500 ;
      RECT 0.0000 381.9500 524.2000 383.0500 ;
      RECT 0.6200 381.6500 524.2000 381.9500 ;
      RECT 0.0000 380.7500 524.2000 381.6500 ;
      RECT 0.0000 380.4500 523.5800 380.7500 ;
      RECT 0.0000 378.1500 524.2000 380.4500 ;
      RECT 0.0000 377.9500 523.5800 378.1500 ;
      RECT 0.6200 377.8500 523.5800 377.9500 ;
      RECT 0.6200 377.6500 524.2000 377.8500 ;
      RECT 0.0000 375.5500 524.2000 377.6500 ;
      RECT 0.0000 375.2500 523.5800 375.5500 ;
      RECT 0.0000 373.9500 524.2000 375.2500 ;
      RECT 0.6200 373.6500 524.2000 373.9500 ;
      RECT 0.0000 372.9500 524.2000 373.6500 ;
      RECT 0.0000 372.6500 523.5800 372.9500 ;
      RECT 0.0000 370.3500 524.2000 372.6500 ;
      RECT 0.0000 370.0500 523.5800 370.3500 ;
      RECT 0.0000 369.9500 524.2000 370.0500 ;
      RECT 0.6200 369.6500 524.2000 369.9500 ;
      RECT 0.0000 367.7500 524.2000 369.6500 ;
      RECT 0.0000 367.4500 523.5800 367.7500 ;
      RECT 0.0000 365.9500 524.2000 367.4500 ;
      RECT 0.6200 365.6500 524.2000 365.9500 ;
      RECT 0.0000 365.1500 524.2000 365.6500 ;
      RECT 0.0000 364.8500 523.5800 365.1500 ;
      RECT 0.0000 362.5500 524.2000 364.8500 ;
      RECT 0.0000 362.2500 523.5800 362.5500 ;
      RECT 0.0000 361.9500 524.2000 362.2500 ;
      RECT 0.6200 361.6500 524.2000 361.9500 ;
      RECT 0.0000 359.9500 524.2000 361.6500 ;
      RECT 0.0000 359.6500 523.5800 359.9500 ;
      RECT 0.0000 357.9500 524.2000 359.6500 ;
      RECT 0.6200 357.6500 524.2000 357.9500 ;
      RECT 0.0000 357.3500 524.2000 357.6500 ;
      RECT 0.0000 357.0500 523.5800 357.3500 ;
      RECT 0.0000 354.7500 524.2000 357.0500 ;
      RECT 0.0000 354.4500 523.5800 354.7500 ;
      RECT 0.0000 353.9500 524.2000 354.4500 ;
      RECT 0.6200 353.6500 524.2000 353.9500 ;
      RECT 0.0000 352.1500 524.2000 353.6500 ;
      RECT 0.0000 351.8500 523.5800 352.1500 ;
      RECT 0.0000 349.9500 524.2000 351.8500 ;
      RECT 0.6200 349.6500 524.2000 349.9500 ;
      RECT 0.0000 349.5500 524.2000 349.6500 ;
      RECT 0.0000 349.2500 523.5800 349.5500 ;
      RECT 0.0000 346.9500 524.2000 349.2500 ;
      RECT 0.0000 346.6500 523.5800 346.9500 ;
      RECT 0.0000 345.9500 524.2000 346.6500 ;
      RECT 0.6200 345.6500 524.2000 345.9500 ;
      RECT 0.0000 344.3500 524.2000 345.6500 ;
      RECT 0.0000 344.0500 523.5800 344.3500 ;
      RECT 0.0000 341.9500 524.2000 344.0500 ;
      RECT 0.6200 341.7500 524.2000 341.9500 ;
      RECT 0.6200 341.6500 523.5800 341.7500 ;
      RECT 0.0000 341.4500 523.5800 341.6500 ;
      RECT 0.0000 339.1500 524.2000 341.4500 ;
      RECT 0.0000 338.8500 523.5800 339.1500 ;
      RECT 0.0000 337.9500 524.2000 338.8500 ;
      RECT 0.6200 337.6500 524.2000 337.9500 ;
      RECT 0.0000 336.5500 524.2000 337.6500 ;
      RECT 0.0000 336.2500 523.5800 336.5500 ;
      RECT 0.0000 333.9500 524.2000 336.2500 ;
      RECT 0.6200 333.6500 523.5800 333.9500 ;
      RECT 0.0000 331.3500 524.2000 333.6500 ;
      RECT 0.0000 331.0500 523.5800 331.3500 ;
      RECT 0.0000 329.9500 524.2000 331.0500 ;
      RECT 0.6200 329.6500 524.2000 329.9500 ;
      RECT 0.0000 328.7500 524.2000 329.6500 ;
      RECT 0.0000 328.4500 523.5800 328.7500 ;
      RECT 0.0000 326.1500 524.2000 328.4500 ;
      RECT 0.0000 325.9500 523.5800 326.1500 ;
      RECT 0.6200 325.8500 523.5800 325.9500 ;
      RECT 0.6200 325.6500 524.2000 325.8500 ;
      RECT 0.0000 323.5500 524.2000 325.6500 ;
      RECT 0.0000 323.2500 523.5800 323.5500 ;
      RECT 0.0000 321.9500 524.2000 323.2500 ;
      RECT 0.6200 321.6500 524.2000 321.9500 ;
      RECT 0.0000 320.9500 524.2000 321.6500 ;
      RECT 0.0000 320.6500 523.5800 320.9500 ;
      RECT 0.0000 318.3500 524.2000 320.6500 ;
      RECT 0.0000 318.0500 523.5800 318.3500 ;
      RECT 0.0000 317.9500 524.2000 318.0500 ;
      RECT 0.6200 317.6500 524.2000 317.9500 ;
      RECT 0.0000 315.7500 524.2000 317.6500 ;
      RECT 0.0000 315.4500 523.5800 315.7500 ;
      RECT 0.0000 313.9500 524.2000 315.4500 ;
      RECT 0.6200 313.6500 524.2000 313.9500 ;
      RECT 0.0000 313.1500 524.2000 313.6500 ;
      RECT 0.0000 312.8500 523.5800 313.1500 ;
      RECT 0.0000 310.5500 524.2000 312.8500 ;
      RECT 0.0000 310.2500 523.5800 310.5500 ;
      RECT 0.0000 309.9500 524.2000 310.2500 ;
      RECT 0.6200 309.6500 524.2000 309.9500 ;
      RECT 0.0000 307.9500 524.2000 309.6500 ;
      RECT 0.0000 307.6500 523.5800 307.9500 ;
      RECT 0.0000 305.9500 524.2000 307.6500 ;
      RECT 0.6200 305.6500 524.2000 305.9500 ;
      RECT 0.0000 305.3500 524.2000 305.6500 ;
      RECT 0.0000 305.0500 523.5800 305.3500 ;
      RECT 0.0000 302.7500 524.2000 305.0500 ;
      RECT 0.0000 302.4500 523.5800 302.7500 ;
      RECT 0.0000 301.9500 524.2000 302.4500 ;
      RECT 0.6200 301.6500 524.2000 301.9500 ;
      RECT 0.0000 300.1500 524.2000 301.6500 ;
      RECT 0.0000 299.8500 523.5800 300.1500 ;
      RECT 0.0000 297.9500 524.2000 299.8500 ;
      RECT 0.6200 297.6500 524.2000 297.9500 ;
      RECT 0.0000 297.5500 524.2000 297.6500 ;
      RECT 0.0000 297.2500 523.5800 297.5500 ;
      RECT 0.0000 294.9500 524.2000 297.2500 ;
      RECT 0.0000 294.6500 523.5800 294.9500 ;
      RECT 0.0000 293.9500 524.2000 294.6500 ;
      RECT 0.6200 293.6500 524.2000 293.9500 ;
      RECT 0.0000 292.3500 524.2000 293.6500 ;
      RECT 0.0000 292.0500 523.5800 292.3500 ;
      RECT 0.0000 289.9500 524.2000 292.0500 ;
      RECT 0.6200 289.7500 524.2000 289.9500 ;
      RECT 0.6200 289.6500 523.5800 289.7500 ;
      RECT 0.0000 289.4500 523.5800 289.6500 ;
      RECT 0.0000 287.1500 524.2000 289.4500 ;
      RECT 0.0000 286.8500 523.5800 287.1500 ;
      RECT 0.0000 285.9500 524.2000 286.8500 ;
      RECT 0.6200 285.6500 524.2000 285.9500 ;
      RECT 0.0000 284.5500 524.2000 285.6500 ;
      RECT 0.0000 284.2500 523.5800 284.5500 ;
      RECT 0.0000 281.9500 524.2000 284.2500 ;
      RECT 0.6200 281.6500 523.5800 281.9500 ;
      RECT 0.0000 279.3500 524.2000 281.6500 ;
      RECT 0.0000 279.0500 523.5800 279.3500 ;
      RECT 0.0000 277.9500 524.2000 279.0500 ;
      RECT 0.6200 277.6500 524.2000 277.9500 ;
      RECT 0.0000 276.7500 524.2000 277.6500 ;
      RECT 0.0000 276.4500 523.5800 276.7500 ;
      RECT 0.0000 274.1500 524.2000 276.4500 ;
      RECT 0.0000 273.9500 523.5800 274.1500 ;
      RECT 0.6200 273.8500 523.5800 273.9500 ;
      RECT 0.6200 273.6500 524.2000 273.8500 ;
      RECT 0.0000 271.5500 524.2000 273.6500 ;
      RECT 0.0000 271.2500 523.5800 271.5500 ;
      RECT 0.0000 269.9500 524.2000 271.2500 ;
      RECT 0.6200 269.6500 524.2000 269.9500 ;
      RECT 0.0000 268.9500 524.2000 269.6500 ;
      RECT 0.0000 268.6500 523.5800 268.9500 ;
      RECT 0.0000 266.3500 524.2000 268.6500 ;
      RECT 0.0000 266.0500 523.5800 266.3500 ;
      RECT 0.0000 265.9500 524.2000 266.0500 ;
      RECT 0.6200 265.6500 524.2000 265.9500 ;
      RECT 0.0000 263.7500 524.2000 265.6500 ;
      RECT 0.0000 263.4500 523.5800 263.7500 ;
      RECT 0.0000 261.9500 524.2000 263.4500 ;
      RECT 0.6200 261.6500 524.2000 261.9500 ;
      RECT 0.0000 261.1500 524.2000 261.6500 ;
      RECT 0.0000 260.8500 523.5800 261.1500 ;
      RECT 0.0000 258.5500 524.2000 260.8500 ;
      RECT 0.0000 258.2500 523.5800 258.5500 ;
      RECT 0.0000 257.9500 524.2000 258.2500 ;
      RECT 0.6200 257.6500 524.2000 257.9500 ;
      RECT 0.0000 255.9500 524.2000 257.6500 ;
      RECT 0.0000 255.6500 523.5800 255.9500 ;
      RECT 0.0000 253.9500 524.2000 255.6500 ;
      RECT 0.6200 253.6500 524.2000 253.9500 ;
      RECT 0.0000 253.3500 524.2000 253.6500 ;
      RECT 0.0000 253.0500 523.5800 253.3500 ;
      RECT 0.0000 250.7500 524.2000 253.0500 ;
      RECT 0.0000 250.4500 523.5800 250.7500 ;
      RECT 0.0000 249.9500 524.2000 250.4500 ;
      RECT 0.6200 249.6500 524.2000 249.9500 ;
      RECT 0.0000 248.1500 524.2000 249.6500 ;
      RECT 0.0000 247.8500 523.5800 248.1500 ;
      RECT 0.0000 245.9500 524.2000 247.8500 ;
      RECT 0.6200 245.6500 524.2000 245.9500 ;
      RECT 0.0000 245.5500 524.2000 245.6500 ;
      RECT 0.0000 245.2500 523.5800 245.5500 ;
      RECT 0.0000 242.9500 524.2000 245.2500 ;
      RECT 0.0000 242.6500 523.5800 242.9500 ;
      RECT 0.0000 241.9500 524.2000 242.6500 ;
      RECT 0.6200 241.6500 524.2000 241.9500 ;
      RECT 0.0000 240.3500 524.2000 241.6500 ;
      RECT 0.0000 240.0500 523.5800 240.3500 ;
      RECT 0.0000 237.9500 524.2000 240.0500 ;
      RECT 0.6200 237.7500 524.2000 237.9500 ;
      RECT 0.6200 237.6500 523.5800 237.7500 ;
      RECT 0.0000 237.4500 523.5800 237.6500 ;
      RECT 0.0000 235.1500 524.2000 237.4500 ;
      RECT 0.0000 234.8500 523.5800 235.1500 ;
      RECT 0.0000 233.9500 524.2000 234.8500 ;
      RECT 0.6200 233.6500 524.2000 233.9500 ;
      RECT 0.0000 232.5500 524.2000 233.6500 ;
      RECT 0.0000 232.2500 523.5800 232.5500 ;
      RECT 0.0000 229.9500 524.2000 232.2500 ;
      RECT 0.6200 229.6500 523.5800 229.9500 ;
      RECT 0.0000 227.3500 524.2000 229.6500 ;
      RECT 0.0000 227.0500 523.5800 227.3500 ;
      RECT 0.0000 225.9500 524.2000 227.0500 ;
      RECT 0.6200 225.6500 524.2000 225.9500 ;
      RECT 0.0000 224.7500 524.2000 225.6500 ;
      RECT 0.0000 224.4500 523.5800 224.7500 ;
      RECT 0.0000 222.1500 524.2000 224.4500 ;
      RECT 0.0000 221.9500 523.5800 222.1500 ;
      RECT 0.6200 221.8500 523.5800 221.9500 ;
      RECT 0.6200 221.6500 524.2000 221.8500 ;
      RECT 0.0000 219.5500 524.2000 221.6500 ;
      RECT 0.0000 219.2500 523.5800 219.5500 ;
      RECT 0.0000 217.9500 524.2000 219.2500 ;
      RECT 0.6200 217.6500 524.2000 217.9500 ;
      RECT 0.0000 216.9500 524.2000 217.6500 ;
      RECT 0.0000 216.6500 523.5800 216.9500 ;
      RECT 0.0000 214.3500 524.2000 216.6500 ;
      RECT 0.0000 214.0500 523.5800 214.3500 ;
      RECT 0.0000 213.9500 524.2000 214.0500 ;
      RECT 0.6200 213.6500 524.2000 213.9500 ;
      RECT 0.0000 211.7500 524.2000 213.6500 ;
      RECT 0.0000 211.4500 523.5800 211.7500 ;
      RECT 0.0000 209.9500 524.2000 211.4500 ;
      RECT 0.6200 209.6500 524.2000 209.9500 ;
      RECT 0.0000 209.1500 524.2000 209.6500 ;
      RECT 0.0000 208.8500 523.5800 209.1500 ;
      RECT 0.0000 206.5500 524.2000 208.8500 ;
      RECT 0.0000 206.2500 523.5800 206.5500 ;
      RECT 0.0000 205.9500 524.2000 206.2500 ;
      RECT 0.6200 205.6500 524.2000 205.9500 ;
      RECT 0.0000 203.9500 524.2000 205.6500 ;
      RECT 0.0000 203.6500 523.5800 203.9500 ;
      RECT 0.0000 201.9500 524.2000 203.6500 ;
      RECT 0.6200 201.6500 524.2000 201.9500 ;
      RECT 0.0000 201.3500 524.2000 201.6500 ;
      RECT 0.0000 201.0500 523.5800 201.3500 ;
      RECT 0.0000 198.7500 524.2000 201.0500 ;
      RECT 0.0000 198.4500 523.5800 198.7500 ;
      RECT 0.0000 197.9500 524.2000 198.4500 ;
      RECT 0.6200 197.6500 524.2000 197.9500 ;
      RECT 0.0000 196.1500 524.2000 197.6500 ;
      RECT 0.0000 195.8500 523.5800 196.1500 ;
      RECT 0.0000 193.9500 524.2000 195.8500 ;
      RECT 0.6200 193.6500 524.2000 193.9500 ;
      RECT 0.0000 193.5500 524.2000 193.6500 ;
      RECT 0.0000 193.2500 523.5800 193.5500 ;
      RECT 0.0000 190.9500 524.2000 193.2500 ;
      RECT 0.0000 190.6500 523.5800 190.9500 ;
      RECT 0.0000 189.9500 524.2000 190.6500 ;
      RECT 0.6200 189.6500 524.2000 189.9500 ;
      RECT 0.0000 188.3500 524.2000 189.6500 ;
      RECT 0.0000 188.0500 523.5800 188.3500 ;
      RECT 0.0000 185.9500 524.2000 188.0500 ;
      RECT 0.6200 185.7500 524.2000 185.9500 ;
      RECT 0.6200 185.6500 523.5800 185.7500 ;
      RECT 0.0000 185.4500 523.5800 185.6500 ;
      RECT 0.0000 183.1500 524.2000 185.4500 ;
      RECT 0.0000 182.8500 523.5800 183.1500 ;
      RECT 0.0000 181.9500 524.2000 182.8500 ;
      RECT 0.6200 181.6500 524.2000 181.9500 ;
      RECT 0.0000 180.5500 524.2000 181.6500 ;
      RECT 0.0000 180.2500 523.5800 180.5500 ;
      RECT 0.0000 177.9500 524.2000 180.2500 ;
      RECT 0.6200 177.6500 523.5800 177.9500 ;
      RECT 0.0000 175.3500 524.2000 177.6500 ;
      RECT 0.0000 175.0500 523.5800 175.3500 ;
      RECT 0.0000 173.9500 524.2000 175.0500 ;
      RECT 0.6200 173.6500 524.2000 173.9500 ;
      RECT 0.0000 172.7500 524.2000 173.6500 ;
      RECT 0.0000 172.4500 523.5800 172.7500 ;
      RECT 0.0000 170.1500 524.2000 172.4500 ;
      RECT 0.0000 169.9500 523.5800 170.1500 ;
      RECT 0.6200 169.8500 523.5800 169.9500 ;
      RECT 0.6200 169.6500 524.2000 169.8500 ;
      RECT 0.0000 167.5500 524.2000 169.6500 ;
      RECT 0.0000 167.2500 523.5800 167.5500 ;
      RECT 0.0000 165.9500 524.2000 167.2500 ;
      RECT 0.6200 165.6500 524.2000 165.9500 ;
      RECT 0.0000 164.9500 524.2000 165.6500 ;
      RECT 0.0000 164.6500 523.5800 164.9500 ;
      RECT 0.0000 162.3500 524.2000 164.6500 ;
      RECT 0.0000 162.0500 523.5800 162.3500 ;
      RECT 0.0000 161.9500 524.2000 162.0500 ;
      RECT 0.6200 161.6500 524.2000 161.9500 ;
      RECT 0.0000 159.7500 524.2000 161.6500 ;
      RECT 0.0000 159.4500 523.5800 159.7500 ;
      RECT 0.0000 157.9500 524.2000 159.4500 ;
      RECT 0.6200 157.6500 524.2000 157.9500 ;
      RECT 0.0000 157.1500 524.2000 157.6500 ;
      RECT 0.0000 156.8500 523.5800 157.1500 ;
      RECT 0.0000 154.5500 524.2000 156.8500 ;
      RECT 0.0000 154.2500 523.5800 154.5500 ;
      RECT 0.0000 153.9500 524.2000 154.2500 ;
      RECT 0.6200 153.6500 524.2000 153.9500 ;
      RECT 0.0000 151.9500 524.2000 153.6500 ;
      RECT 0.0000 151.6500 523.5800 151.9500 ;
      RECT 0.0000 149.9500 524.2000 151.6500 ;
      RECT 0.6200 149.6500 524.2000 149.9500 ;
      RECT 0.0000 149.3500 524.2000 149.6500 ;
      RECT 0.0000 149.0500 523.5800 149.3500 ;
      RECT 0.0000 146.7500 524.2000 149.0500 ;
      RECT 0.0000 146.4500 523.5800 146.7500 ;
      RECT 0.0000 145.9500 524.2000 146.4500 ;
      RECT 0.6200 145.6500 524.2000 145.9500 ;
      RECT 0.0000 144.1500 524.2000 145.6500 ;
      RECT 0.0000 143.8500 523.5800 144.1500 ;
      RECT 0.0000 141.9500 524.2000 143.8500 ;
      RECT 0.6200 141.6500 524.2000 141.9500 ;
      RECT 0.0000 141.5500 524.2000 141.6500 ;
      RECT 0.0000 141.2500 523.5800 141.5500 ;
      RECT 0.0000 138.9500 524.2000 141.2500 ;
      RECT 0.0000 138.6500 523.5800 138.9500 ;
      RECT 0.0000 137.9500 524.2000 138.6500 ;
      RECT 0.6200 137.6500 524.2000 137.9500 ;
      RECT 0.0000 136.3500 524.2000 137.6500 ;
      RECT 0.0000 136.0500 523.5800 136.3500 ;
      RECT 0.0000 133.9500 524.2000 136.0500 ;
      RECT 0.6200 133.7500 524.2000 133.9500 ;
      RECT 0.6200 133.6500 523.5800 133.7500 ;
      RECT 0.0000 133.4500 523.5800 133.6500 ;
      RECT 0.0000 131.1500 524.2000 133.4500 ;
      RECT 0.0000 130.8500 523.5800 131.1500 ;
      RECT 0.0000 129.9500 524.2000 130.8500 ;
      RECT 0.6200 129.6500 524.2000 129.9500 ;
      RECT 0.0000 128.5500 524.2000 129.6500 ;
      RECT 0.0000 128.2500 523.5800 128.5500 ;
      RECT 0.0000 125.9500 524.2000 128.2500 ;
      RECT 0.6200 125.6500 523.5800 125.9500 ;
      RECT 0.0000 123.3500 524.2000 125.6500 ;
      RECT 0.0000 123.0500 523.5800 123.3500 ;
      RECT 0.0000 121.9500 524.2000 123.0500 ;
      RECT 0.6200 121.6500 524.2000 121.9500 ;
      RECT 0.0000 120.7500 524.2000 121.6500 ;
      RECT 0.0000 120.4500 523.5800 120.7500 ;
      RECT 0.0000 118.1500 524.2000 120.4500 ;
      RECT 0.0000 117.9500 523.5800 118.1500 ;
      RECT 0.6200 117.8500 523.5800 117.9500 ;
      RECT 0.6200 117.6500 524.2000 117.8500 ;
      RECT 0.0000 115.5500 524.2000 117.6500 ;
      RECT 0.0000 115.2500 523.5800 115.5500 ;
      RECT 0.0000 113.9500 524.2000 115.2500 ;
      RECT 0.6200 113.6500 524.2000 113.9500 ;
      RECT 0.0000 112.9500 524.2000 113.6500 ;
      RECT 0.0000 112.6500 523.5800 112.9500 ;
      RECT 0.0000 110.3500 524.2000 112.6500 ;
      RECT 0.0000 110.0500 523.5800 110.3500 ;
      RECT 0.0000 109.9500 524.2000 110.0500 ;
      RECT 0.6200 109.6500 524.2000 109.9500 ;
      RECT 0.0000 107.7500 524.2000 109.6500 ;
      RECT 0.0000 107.4500 523.5800 107.7500 ;
      RECT 0.0000 105.9500 524.2000 107.4500 ;
      RECT 0.6200 105.6500 524.2000 105.9500 ;
      RECT 0.0000 105.1500 524.2000 105.6500 ;
      RECT 0.0000 104.8500 523.5800 105.1500 ;
      RECT 0.0000 102.5500 524.2000 104.8500 ;
      RECT 0.0000 102.2500 523.5800 102.5500 ;
      RECT 0.0000 101.9500 524.2000 102.2500 ;
      RECT 0.6200 101.6500 524.2000 101.9500 ;
      RECT 0.0000 99.9500 524.2000 101.6500 ;
      RECT 0.0000 99.6500 523.5800 99.9500 ;
      RECT 0.0000 97.9500 524.2000 99.6500 ;
      RECT 0.6200 97.6500 524.2000 97.9500 ;
      RECT 0.0000 97.3500 524.2000 97.6500 ;
      RECT 0.0000 97.0500 523.5800 97.3500 ;
      RECT 0.0000 94.7500 524.2000 97.0500 ;
      RECT 0.0000 94.4500 523.5800 94.7500 ;
      RECT 0.0000 92.1500 524.2000 94.4500 ;
      RECT 0.0000 91.8500 523.5800 92.1500 ;
      RECT 0.0000 89.5500 524.2000 91.8500 ;
      RECT 0.0000 89.2500 523.5800 89.5500 ;
      RECT 0.0000 86.9500 524.2000 89.2500 ;
      RECT 0.0000 86.6500 523.5800 86.9500 ;
      RECT 0.0000 84.3500 524.2000 86.6500 ;
      RECT 0.0000 84.0500 523.5800 84.3500 ;
      RECT 0.0000 81.7500 524.2000 84.0500 ;
      RECT 0.0000 81.4500 523.5800 81.7500 ;
      RECT 0.0000 79.1500 524.2000 81.4500 ;
      RECT 0.0000 78.8500 523.5800 79.1500 ;
      RECT 0.0000 76.5500 524.2000 78.8500 ;
      RECT 0.0000 76.2500 523.5800 76.5500 ;
      RECT 0.0000 73.9500 524.2000 76.2500 ;
      RECT 0.0000 73.6500 523.5800 73.9500 ;
      RECT 0.0000 71.3500 524.2000 73.6500 ;
      RECT 0.0000 71.0500 523.5800 71.3500 ;
      RECT 0.0000 68.7500 524.2000 71.0500 ;
      RECT 0.0000 68.4500 523.5800 68.7500 ;
      RECT 0.0000 66.1500 524.2000 68.4500 ;
      RECT 0.0000 65.8500 523.5800 66.1500 ;
      RECT 0.0000 63.5500 524.2000 65.8500 ;
      RECT 0.0000 63.2500 523.5800 63.5500 ;
      RECT 0.0000 60.9500 524.2000 63.2500 ;
      RECT 0.0000 60.6500 523.5800 60.9500 ;
      RECT 0.0000 58.3500 524.2000 60.6500 ;
      RECT 0.0000 58.0500 523.5800 58.3500 ;
      RECT 0.0000 55.7500 524.2000 58.0500 ;
      RECT 0.0000 55.4500 523.5800 55.7500 ;
      RECT 0.0000 53.1500 524.2000 55.4500 ;
      RECT 0.0000 52.8500 523.5800 53.1500 ;
      RECT 0.0000 50.5500 524.2000 52.8500 ;
      RECT 0.0000 50.2500 523.5800 50.5500 ;
      RECT 0.0000 47.9500 524.2000 50.2500 ;
      RECT 0.0000 47.6500 523.5800 47.9500 ;
      RECT 0.0000 45.3500 524.2000 47.6500 ;
      RECT 0.0000 45.0500 523.5800 45.3500 ;
      RECT 0.0000 42.7500 524.2000 45.0500 ;
      RECT 0.0000 42.4500 523.5800 42.7500 ;
      RECT 0.0000 40.1500 524.2000 42.4500 ;
      RECT 0.0000 39.8500 523.5800 40.1500 ;
      RECT 0.0000 37.5500 524.2000 39.8500 ;
      RECT 0.0000 37.2500 523.5800 37.5500 ;
      RECT 0.0000 34.9500 524.2000 37.2500 ;
      RECT 0.0000 34.6500 523.5800 34.9500 ;
      RECT 0.0000 32.3500 524.2000 34.6500 ;
      RECT 0.0000 32.0500 523.5800 32.3500 ;
      RECT 0.0000 29.7500 524.2000 32.0500 ;
      RECT 0.0000 29.4500 523.5800 29.7500 ;
      RECT 0.0000 27.1500 524.2000 29.4500 ;
      RECT 0.0000 26.8500 523.5800 27.1500 ;
      RECT 0.0000 24.5500 524.2000 26.8500 ;
      RECT 0.0000 24.2500 523.5800 24.5500 ;
      RECT 0.0000 0.0000 524.2000 24.2500 ;
    LAYER M4 ;
      RECT 0.0000 0.0000 524.2000 524.0000 ;
    LAYER M5 ;
      RECT 0.0000 0.0000 524.2000 524.0000 ;
    LAYER M6 ;
      RECT 0.0000 0.0000 524.2000 524.0000 ;
    LAYER M7 ;
      RECT 0.0000 0.0000 524.2000 524.0000 ;
    LAYER M8 ;
      RECT 0.0000 0.0000 524.2000 524.0000 ;
  END
END core

END LIBRARY
