##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Mon Mar 10 19:44:47 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO sram_w16
  CLASS BLOCK ;
  SIZE 239.8000 BY 239.6000 ;
  FOREIGN sram_w16 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN CLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 69.9500 0.8000 70.0500 ;
    END
  END CLK
  PIN D[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.2500 0.0000 218.3500 0.8000 ;
    END
  END D[127]
  PIN D[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.6500 0.0000 216.7500 0.8000 ;
    END
  END D[126]
  PIN D[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.0500 0.0000 215.1500 0.8000 ;
    END
  END D[125]
  PIN D[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.4500 0.0000 213.5500 0.8000 ;
    END
  END D[124]
  PIN D[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.8500 0.0000 211.9500 0.8000 ;
    END
  END D[123]
  PIN D[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.2500 0.0000 210.3500 0.8000 ;
    END
  END D[122]
  PIN D[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.6500 0.0000 208.7500 0.8000 ;
    END
  END D[121]
  PIN D[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.0500 0.0000 207.1500 0.8000 ;
    END
  END D[120]
  PIN D[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.4500 0.0000 205.5500 0.8000 ;
    END
  END D[119]
  PIN D[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.8500 0.0000 203.9500 0.8000 ;
    END
  END D[118]
  PIN D[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.2500 0.0000 202.3500 0.8000 ;
    END
  END D[117]
  PIN D[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.6500 0.0000 200.7500 0.8000 ;
    END
  END D[116]
  PIN D[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.0500 0.0000 199.1500 0.8000 ;
    END
  END D[115]
  PIN D[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.4500 0.0000 197.5500 0.8000 ;
    END
  END D[114]
  PIN D[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.8500 0.0000 195.9500 0.8000 ;
    END
  END D[113]
  PIN D[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.2500 0.0000 194.3500 0.8000 ;
    END
  END D[112]
  PIN D[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.6500 0.0000 192.7500 0.8000 ;
    END
  END D[111]
  PIN D[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.0500 0.0000 191.1500 0.8000 ;
    END
  END D[110]
  PIN D[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.4500 0.0000 189.5500 0.8000 ;
    END
  END D[109]
  PIN D[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.8500 0.0000 187.9500 0.8000 ;
    END
  END D[108]
  PIN D[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.2500 0.0000 186.3500 0.8000 ;
    END
  END D[107]
  PIN D[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.6500 0.0000 184.7500 0.8000 ;
    END
  END D[106]
  PIN D[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.0500 0.0000 183.1500 0.8000 ;
    END
  END D[105]
  PIN D[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.4500 0.0000 181.5500 0.8000 ;
    END
  END D[104]
  PIN D[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.8500 0.0000 179.9500 0.8000 ;
    END
  END D[103]
  PIN D[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.2500 0.0000 178.3500 0.8000 ;
    END
  END D[102]
  PIN D[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.6500 0.0000 176.7500 0.8000 ;
    END
  END D[101]
  PIN D[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.0500 0.0000 175.1500 0.8000 ;
    END
  END D[100]
  PIN D[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.4500 0.0000 173.5500 0.8000 ;
    END
  END D[99]
  PIN D[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.8500 0.0000 171.9500 0.8000 ;
    END
  END D[98]
  PIN D[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.2500 0.0000 170.3500 0.8000 ;
    END
  END D[97]
  PIN D[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.6500 0.0000 168.7500 0.8000 ;
    END
  END D[96]
  PIN D[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.0500 0.0000 167.1500 0.8000 ;
    END
  END D[95]
  PIN D[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.4500 0.0000 165.5500 0.8000 ;
    END
  END D[94]
  PIN D[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.8500 0.0000 163.9500 0.8000 ;
    END
  END D[93]
  PIN D[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.2500 0.0000 162.3500 0.8000 ;
    END
  END D[92]
  PIN D[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.6500 0.0000 160.7500 0.8000 ;
    END
  END D[91]
  PIN D[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.0500 0.0000 159.1500 0.8000 ;
    END
  END D[90]
  PIN D[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.4500 0.0000 157.5500 0.8000 ;
    END
  END D[89]
  PIN D[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.8500 0.0000 155.9500 0.8000 ;
    END
  END D[88]
  PIN D[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.2500 0.0000 154.3500 0.8000 ;
    END
  END D[87]
  PIN D[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.6500 0.0000 152.7500 0.8000 ;
    END
  END D[86]
  PIN D[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.0500 0.0000 151.1500 0.8000 ;
    END
  END D[85]
  PIN D[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.4500 0.0000 149.5500 0.8000 ;
    END
  END D[84]
  PIN D[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.8500 0.0000 147.9500 0.8000 ;
    END
  END D[83]
  PIN D[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.2500 0.0000 146.3500 0.8000 ;
    END
  END D[82]
  PIN D[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.6500 0.0000 144.7500 0.8000 ;
    END
  END D[81]
  PIN D[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.0500 0.0000 143.1500 0.8000 ;
    END
  END D[80]
  PIN D[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.4500 0.0000 141.5500 0.8000 ;
    END
  END D[79]
  PIN D[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.8500 0.0000 139.9500 0.8000 ;
    END
  END D[78]
  PIN D[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.2500 0.0000 138.3500 0.8000 ;
    END
  END D[77]
  PIN D[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.6500 0.0000 136.7500 0.8000 ;
    END
  END D[76]
  PIN D[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.0500 0.0000 135.1500 0.8000 ;
    END
  END D[75]
  PIN D[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.4500 0.0000 133.5500 0.8000 ;
    END
  END D[74]
  PIN D[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.8500 0.0000 131.9500 0.8000 ;
    END
  END D[73]
  PIN D[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.2500 0.0000 130.3500 0.8000 ;
    END
  END D[72]
  PIN D[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.6500 0.0000 128.7500 0.8000 ;
    END
  END D[71]
  PIN D[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.0500 0.0000 127.1500 0.8000 ;
    END
  END D[70]
  PIN D[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.4500 0.0000 125.5500 0.8000 ;
    END
  END D[69]
  PIN D[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.8500 0.0000 123.9500 0.8000 ;
    END
  END D[68]
  PIN D[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.2500 0.0000 122.3500 0.8000 ;
    END
  END D[67]
  PIN D[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.6500 0.0000 120.7500 0.8000 ;
    END
  END D[66]
  PIN D[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.0500 0.0000 119.1500 0.8000 ;
    END
  END D[65]
  PIN D[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.4500 0.0000 117.5500 0.8000 ;
    END
  END D[64]
  PIN D[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.8500 0.0000 115.9500 0.8000 ;
    END
  END D[63]
  PIN D[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.2500 0.0000 114.3500 0.8000 ;
    END
  END D[62]
  PIN D[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.6500 0.0000 112.7500 0.8000 ;
    END
  END D[61]
  PIN D[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.0500 0.0000 111.1500 0.8000 ;
    END
  END D[60]
  PIN D[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.4500 0.0000 109.5500 0.8000 ;
    END
  END D[59]
  PIN D[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.8500 0.0000 107.9500 0.8000 ;
    END
  END D[58]
  PIN D[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.2500 0.0000 106.3500 0.8000 ;
    END
  END D[57]
  PIN D[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.6500 0.0000 104.7500 0.8000 ;
    END
  END D[56]
  PIN D[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.0500 0.0000 103.1500 0.8000 ;
    END
  END D[55]
  PIN D[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.4500 0.0000 101.5500 0.8000 ;
    END
  END D[54]
  PIN D[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.8500 0.0000 99.9500 0.8000 ;
    END
  END D[53]
  PIN D[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.2500 0.0000 98.3500 0.8000 ;
    END
  END D[52]
  PIN D[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.6500 0.0000 96.7500 0.8000 ;
    END
  END D[51]
  PIN D[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.0500 0.0000 95.1500 0.8000 ;
    END
  END D[50]
  PIN D[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.4500 0.0000 93.5500 0.8000 ;
    END
  END D[49]
  PIN D[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.8500 0.0000 91.9500 0.8000 ;
    END
  END D[48]
  PIN D[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.2500 0.0000 90.3500 0.8000 ;
    END
  END D[47]
  PIN D[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.6500 0.0000 88.7500 0.8000 ;
    END
  END D[46]
  PIN D[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.0500 0.0000 87.1500 0.8000 ;
    END
  END D[45]
  PIN D[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.4500 0.0000 85.5500 0.8000 ;
    END
  END D[44]
  PIN D[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.8500 0.0000 83.9500 0.8000 ;
    END
  END D[43]
  PIN D[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.2500 0.0000 82.3500 0.8000 ;
    END
  END D[42]
  PIN D[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.6500 0.0000 80.7500 0.8000 ;
    END
  END D[41]
  PIN D[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.0500 0.0000 79.1500 0.8000 ;
    END
  END D[40]
  PIN D[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.4500 0.0000 77.5500 0.8000 ;
    END
  END D[39]
  PIN D[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.8500 0.0000 75.9500 0.8000 ;
    END
  END D[38]
  PIN D[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.2500 0.0000 74.3500 0.8000 ;
    END
  END D[37]
  PIN D[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.6500 0.0000 72.7500 0.8000 ;
    END
  END D[36]
  PIN D[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.0500 0.0000 71.1500 0.8000 ;
    END
  END D[35]
  PIN D[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.4500 0.0000 69.5500 0.8000 ;
    END
  END D[34]
  PIN D[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.8500 0.0000 67.9500 0.8000 ;
    END
  END D[33]
  PIN D[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.2500 0.0000 66.3500 0.8000 ;
    END
  END D[32]
  PIN D[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.6500 0.0000 64.7500 0.8000 ;
    END
  END D[31]
  PIN D[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.0500 0.0000 63.1500 0.8000 ;
    END
  END D[30]
  PIN D[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.4500 0.0000 61.5500 0.8000 ;
    END
  END D[29]
  PIN D[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.8500 0.0000 59.9500 0.8000 ;
    END
  END D[28]
  PIN D[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.2500 0.0000 58.3500 0.8000 ;
    END
  END D[27]
  PIN D[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.6500 0.0000 56.7500 0.8000 ;
    END
  END D[26]
  PIN D[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.0500 0.0000 55.1500 0.8000 ;
    END
  END D[25]
  PIN D[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.4500 0.0000 53.5500 0.8000 ;
    END
  END D[24]
  PIN D[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.8500 0.0000 51.9500 0.8000 ;
    END
  END D[23]
  PIN D[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.2500 0.0000 50.3500 0.8000 ;
    END
  END D[22]
  PIN D[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.6500 0.0000 48.7500 0.8000 ;
    END
  END D[21]
  PIN D[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.0500 0.0000 47.1500 0.8000 ;
    END
  END D[20]
  PIN D[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.4500 0.0000 45.5500 0.8000 ;
    END
  END D[19]
  PIN D[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.8500 0.0000 43.9500 0.8000 ;
    END
  END D[18]
  PIN D[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.2500 0.0000 42.3500 0.8000 ;
    END
  END D[17]
  PIN D[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.6500 0.0000 40.7500 0.8000 ;
    END
  END D[16]
  PIN D[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.0500 0.0000 39.1500 0.8000 ;
    END
  END D[15]
  PIN D[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.4500 0.0000 37.5500 0.8000 ;
    END
  END D[14]
  PIN D[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.8500 0.0000 35.9500 0.8000 ;
    END
  END D[13]
  PIN D[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.2500 0.0000 34.3500 0.8000 ;
    END
  END D[12]
  PIN D[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.6500 0.0000 32.7500 0.8000 ;
    END
  END D[11]
  PIN D[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.0500 0.0000 31.1500 0.8000 ;
    END
  END D[10]
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.4500 0.0000 29.5500 0.8000 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.8500 0.0000 27.9500 0.8000 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.2500 0.0000 26.3500 0.8000 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.6500 0.0000 24.7500 0.8000 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.0500 0.0000 23.1500 0.8000 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.4500 0.0000 21.5500 0.8000 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.8500 0.0000 19.9500 0.8000 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.2500 0.0000 18.3500 0.8000 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.6500 0.0000 16.7500 0.8000 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.0500 0.0000 15.1500 0.8000 ;
    END
  END D[0]
  PIN Q[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 218.2500 238.8000 218.3500 239.6000 ;
    END
  END Q[127]
  PIN Q[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 216.6500 238.8000 216.7500 239.6000 ;
    END
  END Q[126]
  PIN Q[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 215.0500 238.8000 215.1500 239.6000 ;
    END
  END Q[125]
  PIN Q[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 213.4500 238.8000 213.5500 239.6000 ;
    END
  END Q[124]
  PIN Q[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 211.8500 238.8000 211.9500 239.6000 ;
    END
  END Q[123]
  PIN Q[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 210.2500 238.8000 210.3500 239.6000 ;
    END
  END Q[122]
  PIN Q[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 208.6500 238.8000 208.7500 239.6000 ;
    END
  END Q[121]
  PIN Q[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 207.0500 238.8000 207.1500 239.6000 ;
    END
  END Q[120]
  PIN Q[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 205.4500 238.8000 205.5500 239.6000 ;
    END
  END Q[119]
  PIN Q[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 203.8500 238.8000 203.9500 239.6000 ;
    END
  END Q[118]
  PIN Q[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 202.2500 238.8000 202.3500 239.6000 ;
    END
  END Q[117]
  PIN Q[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 200.6500 238.8000 200.7500 239.6000 ;
    END
  END Q[116]
  PIN Q[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 199.0500 238.8000 199.1500 239.6000 ;
    END
  END Q[115]
  PIN Q[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 197.4500 238.8000 197.5500 239.6000 ;
    END
  END Q[114]
  PIN Q[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 195.8500 238.8000 195.9500 239.6000 ;
    END
  END Q[113]
  PIN Q[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.2500 238.8000 194.3500 239.6000 ;
    END
  END Q[112]
  PIN Q[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.6500 238.8000 192.7500 239.6000 ;
    END
  END Q[111]
  PIN Q[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.0500 238.8000 191.1500 239.6000 ;
    END
  END Q[110]
  PIN Q[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 189.4500 238.8000 189.5500 239.6000 ;
    END
  END Q[109]
  PIN Q[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.8500 238.8000 187.9500 239.6000 ;
    END
  END Q[108]
  PIN Q[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 186.2500 238.8000 186.3500 239.6000 ;
    END
  END Q[107]
  PIN Q[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 184.6500 238.8000 184.7500 239.6000 ;
    END
  END Q[106]
  PIN Q[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 183.0500 238.8000 183.1500 239.6000 ;
    END
  END Q[105]
  PIN Q[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.4500 238.8000 181.5500 239.6000 ;
    END
  END Q[104]
  PIN Q[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 179.8500 238.8000 179.9500 239.6000 ;
    END
  END Q[103]
  PIN Q[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.2500 238.8000 178.3500 239.6000 ;
    END
  END Q[102]
  PIN Q[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 176.6500 238.8000 176.7500 239.6000 ;
    END
  END Q[101]
  PIN Q[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 175.0500 238.8000 175.1500 239.6000 ;
    END
  END Q[100]
  PIN Q[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 173.4500 238.8000 173.5500 239.6000 ;
    END
  END Q[99]
  PIN Q[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.8500 238.8000 171.9500 239.6000 ;
    END
  END Q[98]
  PIN Q[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 170.2500 238.8000 170.3500 239.6000 ;
    END
  END Q[97]
  PIN Q[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 168.6500 238.8000 168.7500 239.6000 ;
    END
  END Q[96]
  PIN Q[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.0500 238.8000 167.1500 239.6000 ;
    END
  END Q[95]
  PIN Q[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 165.4500 238.8000 165.5500 239.6000 ;
    END
  END Q[94]
  PIN Q[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 163.8500 238.8000 163.9500 239.6000 ;
    END
  END Q[93]
  PIN Q[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 162.2500 238.8000 162.3500 239.6000 ;
    END
  END Q[92]
  PIN Q[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 160.6500 238.8000 160.7500 239.6000 ;
    END
  END Q[91]
  PIN Q[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 159.0500 238.8000 159.1500 239.6000 ;
    END
  END Q[90]
  PIN Q[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 157.4500 238.8000 157.5500 239.6000 ;
    END
  END Q[89]
  PIN Q[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 155.8500 238.8000 155.9500 239.6000 ;
    END
  END Q[88]
  PIN Q[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 154.2500 238.8000 154.3500 239.6000 ;
    END
  END Q[87]
  PIN Q[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 152.6500 238.8000 152.7500 239.6000 ;
    END
  END Q[86]
  PIN Q[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 151.0500 238.8000 151.1500 239.6000 ;
    END
  END Q[85]
  PIN Q[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 149.4500 238.8000 149.5500 239.6000 ;
    END
  END Q[84]
  PIN Q[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 147.8500 238.8000 147.9500 239.6000 ;
    END
  END Q[83]
  PIN Q[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 146.2500 238.8000 146.3500 239.6000 ;
    END
  END Q[82]
  PIN Q[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 144.6500 238.8000 144.7500 239.6000 ;
    END
  END Q[81]
  PIN Q[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 143.0500 238.8000 143.1500 239.6000 ;
    END
  END Q[80]
  PIN Q[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 141.4500 238.8000 141.5500 239.6000 ;
    END
  END Q[79]
  PIN Q[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 139.8500 238.8000 139.9500 239.6000 ;
    END
  END Q[78]
  PIN Q[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 138.2500 238.8000 138.3500 239.6000 ;
    END
  END Q[77]
  PIN Q[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 136.6500 238.8000 136.7500 239.6000 ;
    END
  END Q[76]
  PIN Q[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 135.0500 238.8000 135.1500 239.6000 ;
    END
  END Q[75]
  PIN Q[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.4500 238.8000 133.5500 239.6000 ;
    END
  END Q[74]
  PIN Q[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 131.8500 238.8000 131.9500 239.6000 ;
    END
  END Q[73]
  PIN Q[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 130.2500 238.8000 130.3500 239.6000 ;
    END
  END Q[72]
  PIN Q[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 128.6500 238.8000 128.7500 239.6000 ;
    END
  END Q[71]
  PIN Q[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.0500 238.8000 127.1500 239.6000 ;
    END
  END Q[70]
  PIN Q[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 125.4500 238.8000 125.5500 239.6000 ;
    END
  END Q[69]
  PIN Q[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.8500 238.8000 123.9500 239.6000 ;
    END
  END Q[68]
  PIN Q[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 122.2500 238.8000 122.3500 239.6000 ;
    END
  END Q[67]
  PIN Q[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 120.6500 238.8000 120.7500 239.6000 ;
    END
  END Q[66]
  PIN Q[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.0500 238.8000 119.1500 239.6000 ;
    END
  END Q[65]
  PIN Q[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 117.4500 238.8000 117.5500 239.6000 ;
    END
  END Q[64]
  PIN Q[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 115.8500 238.8000 115.9500 239.6000 ;
    END
  END Q[63]
  PIN Q[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 114.2500 238.8000 114.3500 239.6000 ;
    END
  END Q[62]
  PIN Q[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 112.6500 238.8000 112.7500 239.6000 ;
    END
  END Q[61]
  PIN Q[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 111.0500 238.8000 111.1500 239.6000 ;
    END
  END Q[60]
  PIN Q[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 109.4500 238.8000 109.5500 239.6000 ;
    END
  END Q[59]
  PIN Q[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 107.8500 238.8000 107.9500 239.6000 ;
    END
  END Q[58]
  PIN Q[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.2500 238.8000 106.3500 239.6000 ;
    END
  END Q[57]
  PIN Q[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.6500 238.8000 104.7500 239.6000 ;
    END
  END Q[56]
  PIN Q[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 103.0500 238.8000 103.1500 239.6000 ;
    END
  END Q[55]
  PIN Q[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 101.4500 238.8000 101.5500 239.6000 ;
    END
  END Q[54]
  PIN Q[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 99.8500 238.8000 99.9500 239.6000 ;
    END
  END Q[53]
  PIN Q[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 98.2500 238.8000 98.3500 239.6000 ;
    END
  END Q[52]
  PIN Q[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 96.6500 238.8000 96.7500 239.6000 ;
    END
  END Q[51]
  PIN Q[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 95.0500 238.8000 95.1500 239.6000 ;
    END
  END Q[50]
  PIN Q[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 93.4500 238.8000 93.5500 239.6000 ;
    END
  END Q[49]
  PIN Q[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 91.8500 238.8000 91.9500 239.6000 ;
    END
  END Q[48]
  PIN Q[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 90.2500 238.8000 90.3500 239.6000 ;
    END
  END Q[47]
  PIN Q[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 88.6500 238.8000 88.7500 239.6000 ;
    END
  END Q[46]
  PIN Q[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 87.0500 238.8000 87.1500 239.6000 ;
    END
  END Q[45]
  PIN Q[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 85.4500 238.8000 85.5500 239.6000 ;
    END
  END Q[44]
  PIN Q[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 83.8500 238.8000 83.9500 239.6000 ;
    END
  END Q[43]
  PIN Q[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 82.2500 238.8000 82.3500 239.6000 ;
    END
  END Q[42]
  PIN Q[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 80.6500 238.8000 80.7500 239.6000 ;
    END
  END Q[41]
  PIN Q[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 79.0500 238.8000 79.1500 239.6000 ;
    END
  END Q[40]
  PIN Q[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.4500 238.8000 77.5500 239.6000 ;
    END
  END Q[39]
  PIN Q[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.8500 238.8000 75.9500 239.6000 ;
    END
  END Q[38]
  PIN Q[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 74.2500 238.8000 74.3500 239.6000 ;
    END
  END Q[37]
  PIN Q[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 72.6500 238.8000 72.7500 239.6000 ;
    END
  END Q[36]
  PIN Q[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 71.0500 238.8000 71.1500 239.6000 ;
    END
  END Q[35]
  PIN Q[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 69.4500 238.8000 69.5500 239.6000 ;
    END
  END Q[34]
  PIN Q[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 67.8500 238.8000 67.9500 239.6000 ;
    END
  END Q[33]
  PIN Q[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 66.2500 238.8000 66.3500 239.6000 ;
    END
  END Q[32]
  PIN Q[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 64.6500 238.8000 64.7500 239.6000 ;
    END
  END Q[31]
  PIN Q[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 63.0500 238.8000 63.1500 239.6000 ;
    END
  END Q[30]
  PIN Q[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 61.4500 238.8000 61.5500 239.6000 ;
    END
  END Q[29]
  PIN Q[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 59.8500 238.8000 59.9500 239.6000 ;
    END
  END Q[28]
  PIN Q[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 58.2500 238.8000 58.3500 239.6000 ;
    END
  END Q[27]
  PIN Q[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 56.6500 238.8000 56.7500 239.6000 ;
    END
  END Q[26]
  PIN Q[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 55.0500 238.8000 55.1500 239.6000 ;
    END
  END Q[25]
  PIN Q[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 53.4500 238.8000 53.5500 239.6000 ;
    END
  END Q[24]
  PIN Q[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 51.8500 238.8000 51.9500 239.6000 ;
    END
  END Q[23]
  PIN Q[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 50.2500 238.8000 50.3500 239.6000 ;
    END
  END Q[22]
  PIN Q[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 48.6500 238.8000 48.7500 239.6000 ;
    END
  END Q[21]
  PIN Q[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 47.0500 238.8000 47.1500 239.6000 ;
    END
  END Q[20]
  PIN Q[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 45.4500 238.8000 45.5500 239.6000 ;
    END
  END Q[19]
  PIN Q[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 43.8500 238.8000 43.9500 239.6000 ;
    END
  END Q[18]
  PIN Q[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 42.2500 238.8000 42.3500 239.6000 ;
    END
  END Q[17]
  PIN Q[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 40.6500 238.8000 40.7500 239.6000 ;
    END
  END Q[16]
  PIN Q[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 39.0500 238.8000 39.1500 239.6000 ;
    END
  END Q[15]
  PIN Q[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 37.4500 238.8000 37.5500 239.6000 ;
    END
  END Q[14]
  PIN Q[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 35.8500 238.8000 35.9500 239.6000 ;
    END
  END Q[13]
  PIN Q[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 34.2500 238.8000 34.3500 239.6000 ;
    END
  END Q[12]
  PIN Q[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 32.6500 238.8000 32.7500 239.6000 ;
    END
  END Q[11]
  PIN Q[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 31.0500 238.8000 31.1500 239.6000 ;
    END
  END Q[10]
  PIN Q[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 29.4500 238.8000 29.5500 239.6000 ;
    END
  END Q[9]
  PIN Q[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 27.8500 238.8000 27.9500 239.6000 ;
    END
  END Q[8]
  PIN Q[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 26.2500 238.8000 26.3500 239.6000 ;
    END
  END Q[7]
  PIN Q[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 24.6500 238.8000 24.7500 239.6000 ;
    END
  END Q[6]
  PIN Q[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 23.0500 238.8000 23.1500 239.6000 ;
    END
  END Q[5]
  PIN Q[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 21.4500 238.8000 21.5500 239.6000 ;
    END
  END Q[4]
  PIN Q[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 19.8500 238.8000 19.9500 239.6000 ;
    END
  END Q[3]
  PIN Q[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 18.2500 238.8000 18.3500 239.6000 ;
    END
  END Q[2]
  PIN Q[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 16.6500 238.8000 16.7500 239.6000 ;
    END
  END Q[1]
  PIN Q[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 15.0500 238.8000 15.1500 239.6000 ;
    END
  END Q[0]
  PIN CEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 65.9500 0.8000 66.0500 ;
    END
  END CEN
  PIN WEN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 73.9500 0.8000 74.0500 ;
    END
  END WEN
  PIN A[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 61.9500 0.8000 62.0500 ;
    END
  END A[3]
  PIN A[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.9500 0.8000 58.0500 ;
    END
  END A[2]
  PIN A[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 53.9500 0.8000 54.0500 ;
    END
  END A[1]
  PIN A[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 49.9500 0.8000 50.0500 ;
    END
  END A[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 28.0000 10.0000 30.0000 229.6000 ;
        RECT 56.0550 10.0000 58.0550 229.6000 ;
        RECT 84.1100 10.0000 86.1100 229.6000 ;
        RECT 112.1650 10.0000 114.1650 229.6000 ;
        RECT 140.2200 10.0000 142.2200 229.6000 ;
        RECT 168.2750 10.0000 170.2750 229.6000 ;
        RECT 196.3300 10.0000 198.3300 229.6000 ;
        RECT 224.3850 10.0000 226.3850 229.6000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 20.0000 10.0000 22.0000 229.6000 ;
        RECT 48.0550 10.0000 50.0550 229.6000 ;
        RECT 76.1100 10.0000 78.1100 229.6000 ;
        RECT 104.1650 10.0000 106.1650 229.6000 ;
        RECT 132.2200 10.0000 134.2200 229.6000 ;
        RECT 160.2750 10.0000 162.2750 229.6000 ;
        RECT 188.3300 10.0000 190.3300 229.6000 ;
        RECT 216.3850 10.0000 218.3850 229.6000 ;
        RECT 20.0000 9.8350 22.0000 10.1650 ;
        RECT 48.0550 9.8350 50.0550 10.1650 ;
        RECT 76.1100 9.8350 78.1100 10.1650 ;
        RECT 104.1650 9.8350 106.1650 10.1650 ;
        RECT 132.2200 9.8350 134.2200 10.1650 ;
        RECT 160.2750 9.8350 162.2750 10.1650 ;
        RECT 188.3300 9.8350 190.3300 10.1650 ;
        RECT 216.3850 9.8350 218.3850 10.1650 ;
        RECT 20.0000 229.4350 22.0000 229.7650 ;
        RECT 48.0550 229.4350 50.0550 229.7650 ;
        RECT 76.1100 229.4350 78.1100 229.7650 ;
        RECT 104.1650 229.4350 106.1650 229.7650 ;
        RECT 132.2200 229.4350 134.2200 229.7650 ;
        RECT 160.2750 229.4350 162.2750 229.7650 ;
        RECT 188.3300 229.4350 190.3300 229.7650 ;
        RECT 216.3850 229.4350 218.3850 229.7650 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 239.8000 239.6000 ;
    LAYER M2 ;
      RECT 218.4500 238.7000 239.8000 239.6000 ;
      RECT 216.8500 238.7000 218.1500 239.6000 ;
      RECT 215.2500 238.7000 216.5500 239.6000 ;
      RECT 213.6500 238.7000 214.9500 239.6000 ;
      RECT 212.0500 238.7000 213.3500 239.6000 ;
      RECT 210.4500 238.7000 211.7500 239.6000 ;
      RECT 208.8500 238.7000 210.1500 239.6000 ;
      RECT 207.2500 238.7000 208.5500 239.6000 ;
      RECT 205.6500 238.7000 206.9500 239.6000 ;
      RECT 204.0500 238.7000 205.3500 239.6000 ;
      RECT 202.4500 238.7000 203.7500 239.6000 ;
      RECT 200.8500 238.7000 202.1500 239.6000 ;
      RECT 199.2500 238.7000 200.5500 239.6000 ;
      RECT 197.6500 238.7000 198.9500 239.6000 ;
      RECT 196.0500 238.7000 197.3500 239.6000 ;
      RECT 194.4500 238.7000 195.7500 239.6000 ;
      RECT 192.8500 238.7000 194.1500 239.6000 ;
      RECT 191.2500 238.7000 192.5500 239.6000 ;
      RECT 189.6500 238.7000 190.9500 239.6000 ;
      RECT 188.0500 238.7000 189.3500 239.6000 ;
      RECT 186.4500 238.7000 187.7500 239.6000 ;
      RECT 184.8500 238.7000 186.1500 239.6000 ;
      RECT 183.2500 238.7000 184.5500 239.6000 ;
      RECT 181.6500 238.7000 182.9500 239.6000 ;
      RECT 180.0500 238.7000 181.3500 239.6000 ;
      RECT 178.4500 238.7000 179.7500 239.6000 ;
      RECT 176.8500 238.7000 178.1500 239.6000 ;
      RECT 175.2500 238.7000 176.5500 239.6000 ;
      RECT 173.6500 238.7000 174.9500 239.6000 ;
      RECT 172.0500 238.7000 173.3500 239.6000 ;
      RECT 170.4500 238.7000 171.7500 239.6000 ;
      RECT 168.8500 238.7000 170.1500 239.6000 ;
      RECT 167.2500 238.7000 168.5500 239.6000 ;
      RECT 165.6500 238.7000 166.9500 239.6000 ;
      RECT 164.0500 238.7000 165.3500 239.6000 ;
      RECT 162.4500 238.7000 163.7500 239.6000 ;
      RECT 160.8500 238.7000 162.1500 239.6000 ;
      RECT 159.2500 238.7000 160.5500 239.6000 ;
      RECT 157.6500 238.7000 158.9500 239.6000 ;
      RECT 156.0500 238.7000 157.3500 239.6000 ;
      RECT 154.4500 238.7000 155.7500 239.6000 ;
      RECT 152.8500 238.7000 154.1500 239.6000 ;
      RECT 151.2500 238.7000 152.5500 239.6000 ;
      RECT 149.6500 238.7000 150.9500 239.6000 ;
      RECT 148.0500 238.7000 149.3500 239.6000 ;
      RECT 146.4500 238.7000 147.7500 239.6000 ;
      RECT 144.8500 238.7000 146.1500 239.6000 ;
      RECT 143.2500 238.7000 144.5500 239.6000 ;
      RECT 141.6500 238.7000 142.9500 239.6000 ;
      RECT 140.0500 238.7000 141.3500 239.6000 ;
      RECT 138.4500 238.7000 139.7500 239.6000 ;
      RECT 136.8500 238.7000 138.1500 239.6000 ;
      RECT 135.2500 238.7000 136.5500 239.6000 ;
      RECT 133.6500 238.7000 134.9500 239.6000 ;
      RECT 132.0500 238.7000 133.3500 239.6000 ;
      RECT 130.4500 238.7000 131.7500 239.6000 ;
      RECT 128.8500 238.7000 130.1500 239.6000 ;
      RECT 127.2500 238.7000 128.5500 239.6000 ;
      RECT 125.6500 238.7000 126.9500 239.6000 ;
      RECT 124.0500 238.7000 125.3500 239.6000 ;
      RECT 122.4500 238.7000 123.7500 239.6000 ;
      RECT 120.8500 238.7000 122.1500 239.6000 ;
      RECT 119.2500 238.7000 120.5500 239.6000 ;
      RECT 117.6500 238.7000 118.9500 239.6000 ;
      RECT 116.0500 238.7000 117.3500 239.6000 ;
      RECT 114.4500 238.7000 115.7500 239.6000 ;
      RECT 112.8500 238.7000 114.1500 239.6000 ;
      RECT 111.2500 238.7000 112.5500 239.6000 ;
      RECT 109.6500 238.7000 110.9500 239.6000 ;
      RECT 108.0500 238.7000 109.3500 239.6000 ;
      RECT 106.4500 238.7000 107.7500 239.6000 ;
      RECT 104.8500 238.7000 106.1500 239.6000 ;
      RECT 103.2500 238.7000 104.5500 239.6000 ;
      RECT 101.6500 238.7000 102.9500 239.6000 ;
      RECT 100.0500 238.7000 101.3500 239.6000 ;
      RECT 98.4500 238.7000 99.7500 239.6000 ;
      RECT 96.8500 238.7000 98.1500 239.6000 ;
      RECT 95.2500 238.7000 96.5500 239.6000 ;
      RECT 93.6500 238.7000 94.9500 239.6000 ;
      RECT 92.0500 238.7000 93.3500 239.6000 ;
      RECT 90.4500 238.7000 91.7500 239.6000 ;
      RECT 88.8500 238.7000 90.1500 239.6000 ;
      RECT 87.2500 238.7000 88.5500 239.6000 ;
      RECT 85.6500 238.7000 86.9500 239.6000 ;
      RECT 84.0500 238.7000 85.3500 239.6000 ;
      RECT 82.4500 238.7000 83.7500 239.6000 ;
      RECT 80.8500 238.7000 82.1500 239.6000 ;
      RECT 79.2500 238.7000 80.5500 239.6000 ;
      RECT 77.6500 238.7000 78.9500 239.6000 ;
      RECT 76.0500 238.7000 77.3500 239.6000 ;
      RECT 74.4500 238.7000 75.7500 239.6000 ;
      RECT 72.8500 238.7000 74.1500 239.6000 ;
      RECT 71.2500 238.7000 72.5500 239.6000 ;
      RECT 69.6500 238.7000 70.9500 239.6000 ;
      RECT 68.0500 238.7000 69.3500 239.6000 ;
      RECT 66.4500 238.7000 67.7500 239.6000 ;
      RECT 64.8500 238.7000 66.1500 239.6000 ;
      RECT 63.2500 238.7000 64.5500 239.6000 ;
      RECT 61.6500 238.7000 62.9500 239.6000 ;
      RECT 60.0500 238.7000 61.3500 239.6000 ;
      RECT 58.4500 238.7000 59.7500 239.6000 ;
      RECT 56.8500 238.7000 58.1500 239.6000 ;
      RECT 55.2500 238.7000 56.5500 239.6000 ;
      RECT 53.6500 238.7000 54.9500 239.6000 ;
      RECT 52.0500 238.7000 53.3500 239.6000 ;
      RECT 50.4500 238.7000 51.7500 239.6000 ;
      RECT 48.8500 238.7000 50.1500 239.6000 ;
      RECT 47.2500 238.7000 48.5500 239.6000 ;
      RECT 45.6500 238.7000 46.9500 239.6000 ;
      RECT 44.0500 238.7000 45.3500 239.6000 ;
      RECT 42.4500 238.7000 43.7500 239.6000 ;
      RECT 40.8500 238.7000 42.1500 239.6000 ;
      RECT 39.2500 238.7000 40.5500 239.6000 ;
      RECT 37.6500 238.7000 38.9500 239.6000 ;
      RECT 36.0500 238.7000 37.3500 239.6000 ;
      RECT 34.4500 238.7000 35.7500 239.6000 ;
      RECT 32.8500 238.7000 34.1500 239.6000 ;
      RECT 31.2500 238.7000 32.5500 239.6000 ;
      RECT 29.6500 238.7000 30.9500 239.6000 ;
      RECT 28.0500 238.7000 29.3500 239.6000 ;
      RECT 26.4500 238.7000 27.7500 239.6000 ;
      RECT 24.8500 238.7000 26.1500 239.6000 ;
      RECT 23.2500 238.7000 24.5500 239.6000 ;
      RECT 21.6500 238.7000 22.9500 239.6000 ;
      RECT 20.0500 238.7000 21.3500 239.6000 ;
      RECT 18.4500 238.7000 19.7500 239.6000 ;
      RECT 16.8500 238.7000 18.1500 239.6000 ;
      RECT 15.2500 238.7000 16.5500 239.6000 ;
      RECT 0.0000 238.7000 14.9500 239.6000 ;
      RECT 0.0000 0.9000 239.8000 238.7000 ;
      RECT 218.4500 0.0000 239.8000 0.9000 ;
      RECT 216.8500 0.0000 218.1500 0.9000 ;
      RECT 215.2500 0.0000 216.5500 0.9000 ;
      RECT 213.6500 0.0000 214.9500 0.9000 ;
      RECT 212.0500 0.0000 213.3500 0.9000 ;
      RECT 210.4500 0.0000 211.7500 0.9000 ;
      RECT 208.8500 0.0000 210.1500 0.9000 ;
      RECT 207.2500 0.0000 208.5500 0.9000 ;
      RECT 205.6500 0.0000 206.9500 0.9000 ;
      RECT 204.0500 0.0000 205.3500 0.9000 ;
      RECT 202.4500 0.0000 203.7500 0.9000 ;
      RECT 200.8500 0.0000 202.1500 0.9000 ;
      RECT 199.2500 0.0000 200.5500 0.9000 ;
      RECT 197.6500 0.0000 198.9500 0.9000 ;
      RECT 196.0500 0.0000 197.3500 0.9000 ;
      RECT 194.4500 0.0000 195.7500 0.9000 ;
      RECT 192.8500 0.0000 194.1500 0.9000 ;
      RECT 191.2500 0.0000 192.5500 0.9000 ;
      RECT 189.6500 0.0000 190.9500 0.9000 ;
      RECT 188.0500 0.0000 189.3500 0.9000 ;
      RECT 186.4500 0.0000 187.7500 0.9000 ;
      RECT 184.8500 0.0000 186.1500 0.9000 ;
      RECT 183.2500 0.0000 184.5500 0.9000 ;
      RECT 181.6500 0.0000 182.9500 0.9000 ;
      RECT 180.0500 0.0000 181.3500 0.9000 ;
      RECT 178.4500 0.0000 179.7500 0.9000 ;
      RECT 176.8500 0.0000 178.1500 0.9000 ;
      RECT 175.2500 0.0000 176.5500 0.9000 ;
      RECT 173.6500 0.0000 174.9500 0.9000 ;
      RECT 172.0500 0.0000 173.3500 0.9000 ;
      RECT 170.4500 0.0000 171.7500 0.9000 ;
      RECT 168.8500 0.0000 170.1500 0.9000 ;
      RECT 167.2500 0.0000 168.5500 0.9000 ;
      RECT 165.6500 0.0000 166.9500 0.9000 ;
      RECT 164.0500 0.0000 165.3500 0.9000 ;
      RECT 162.4500 0.0000 163.7500 0.9000 ;
      RECT 160.8500 0.0000 162.1500 0.9000 ;
      RECT 159.2500 0.0000 160.5500 0.9000 ;
      RECT 157.6500 0.0000 158.9500 0.9000 ;
      RECT 156.0500 0.0000 157.3500 0.9000 ;
      RECT 154.4500 0.0000 155.7500 0.9000 ;
      RECT 152.8500 0.0000 154.1500 0.9000 ;
      RECT 151.2500 0.0000 152.5500 0.9000 ;
      RECT 149.6500 0.0000 150.9500 0.9000 ;
      RECT 148.0500 0.0000 149.3500 0.9000 ;
      RECT 146.4500 0.0000 147.7500 0.9000 ;
      RECT 144.8500 0.0000 146.1500 0.9000 ;
      RECT 143.2500 0.0000 144.5500 0.9000 ;
      RECT 141.6500 0.0000 142.9500 0.9000 ;
      RECT 140.0500 0.0000 141.3500 0.9000 ;
      RECT 138.4500 0.0000 139.7500 0.9000 ;
      RECT 136.8500 0.0000 138.1500 0.9000 ;
      RECT 135.2500 0.0000 136.5500 0.9000 ;
      RECT 133.6500 0.0000 134.9500 0.9000 ;
      RECT 132.0500 0.0000 133.3500 0.9000 ;
      RECT 130.4500 0.0000 131.7500 0.9000 ;
      RECT 128.8500 0.0000 130.1500 0.9000 ;
      RECT 127.2500 0.0000 128.5500 0.9000 ;
      RECT 125.6500 0.0000 126.9500 0.9000 ;
      RECT 124.0500 0.0000 125.3500 0.9000 ;
      RECT 122.4500 0.0000 123.7500 0.9000 ;
      RECT 120.8500 0.0000 122.1500 0.9000 ;
      RECT 119.2500 0.0000 120.5500 0.9000 ;
      RECT 117.6500 0.0000 118.9500 0.9000 ;
      RECT 116.0500 0.0000 117.3500 0.9000 ;
      RECT 114.4500 0.0000 115.7500 0.9000 ;
      RECT 112.8500 0.0000 114.1500 0.9000 ;
      RECT 111.2500 0.0000 112.5500 0.9000 ;
      RECT 109.6500 0.0000 110.9500 0.9000 ;
      RECT 108.0500 0.0000 109.3500 0.9000 ;
      RECT 106.4500 0.0000 107.7500 0.9000 ;
      RECT 104.8500 0.0000 106.1500 0.9000 ;
      RECT 103.2500 0.0000 104.5500 0.9000 ;
      RECT 101.6500 0.0000 102.9500 0.9000 ;
      RECT 100.0500 0.0000 101.3500 0.9000 ;
      RECT 98.4500 0.0000 99.7500 0.9000 ;
      RECT 96.8500 0.0000 98.1500 0.9000 ;
      RECT 95.2500 0.0000 96.5500 0.9000 ;
      RECT 93.6500 0.0000 94.9500 0.9000 ;
      RECT 92.0500 0.0000 93.3500 0.9000 ;
      RECT 90.4500 0.0000 91.7500 0.9000 ;
      RECT 88.8500 0.0000 90.1500 0.9000 ;
      RECT 87.2500 0.0000 88.5500 0.9000 ;
      RECT 85.6500 0.0000 86.9500 0.9000 ;
      RECT 84.0500 0.0000 85.3500 0.9000 ;
      RECT 82.4500 0.0000 83.7500 0.9000 ;
      RECT 80.8500 0.0000 82.1500 0.9000 ;
      RECT 79.2500 0.0000 80.5500 0.9000 ;
      RECT 77.6500 0.0000 78.9500 0.9000 ;
      RECT 76.0500 0.0000 77.3500 0.9000 ;
      RECT 74.4500 0.0000 75.7500 0.9000 ;
      RECT 72.8500 0.0000 74.1500 0.9000 ;
      RECT 71.2500 0.0000 72.5500 0.9000 ;
      RECT 69.6500 0.0000 70.9500 0.9000 ;
      RECT 68.0500 0.0000 69.3500 0.9000 ;
      RECT 66.4500 0.0000 67.7500 0.9000 ;
      RECT 64.8500 0.0000 66.1500 0.9000 ;
      RECT 63.2500 0.0000 64.5500 0.9000 ;
      RECT 61.6500 0.0000 62.9500 0.9000 ;
      RECT 60.0500 0.0000 61.3500 0.9000 ;
      RECT 58.4500 0.0000 59.7500 0.9000 ;
      RECT 56.8500 0.0000 58.1500 0.9000 ;
      RECT 55.2500 0.0000 56.5500 0.9000 ;
      RECT 53.6500 0.0000 54.9500 0.9000 ;
      RECT 52.0500 0.0000 53.3500 0.9000 ;
      RECT 50.4500 0.0000 51.7500 0.9000 ;
      RECT 48.8500 0.0000 50.1500 0.9000 ;
      RECT 47.2500 0.0000 48.5500 0.9000 ;
      RECT 45.6500 0.0000 46.9500 0.9000 ;
      RECT 44.0500 0.0000 45.3500 0.9000 ;
      RECT 42.4500 0.0000 43.7500 0.9000 ;
      RECT 40.8500 0.0000 42.1500 0.9000 ;
      RECT 39.2500 0.0000 40.5500 0.9000 ;
      RECT 37.6500 0.0000 38.9500 0.9000 ;
      RECT 36.0500 0.0000 37.3500 0.9000 ;
      RECT 34.4500 0.0000 35.7500 0.9000 ;
      RECT 32.8500 0.0000 34.1500 0.9000 ;
      RECT 31.2500 0.0000 32.5500 0.9000 ;
      RECT 29.6500 0.0000 30.9500 0.9000 ;
      RECT 28.0500 0.0000 29.3500 0.9000 ;
      RECT 26.4500 0.0000 27.7500 0.9000 ;
      RECT 24.8500 0.0000 26.1500 0.9000 ;
      RECT 23.2500 0.0000 24.5500 0.9000 ;
      RECT 21.6500 0.0000 22.9500 0.9000 ;
      RECT 20.0500 0.0000 21.3500 0.9000 ;
      RECT 18.4500 0.0000 19.7500 0.9000 ;
      RECT 16.8500 0.0000 18.1500 0.9000 ;
      RECT 15.2500 0.0000 16.5500 0.9000 ;
      RECT 0.0000 0.0000 14.9500 0.9000 ;
    LAYER M3 ;
      RECT 0.0000 74.1500 239.8000 239.6000 ;
      RECT 0.9000 73.8500 239.8000 74.1500 ;
      RECT 0.0000 70.1500 239.8000 73.8500 ;
      RECT 0.9000 69.8500 239.8000 70.1500 ;
      RECT 0.0000 66.1500 239.8000 69.8500 ;
      RECT 0.9000 65.8500 239.8000 66.1500 ;
      RECT 0.0000 62.1500 239.8000 65.8500 ;
      RECT 0.9000 61.8500 239.8000 62.1500 ;
      RECT 0.0000 58.1500 239.8000 61.8500 ;
      RECT 0.9000 57.8500 239.8000 58.1500 ;
      RECT 0.0000 54.1500 239.8000 57.8500 ;
      RECT 0.9000 53.8500 239.8000 54.1500 ;
      RECT 0.0000 50.1500 239.8000 53.8500 ;
      RECT 0.9000 49.8500 239.8000 50.1500 ;
      RECT 0.0000 0.0000 239.8000 49.8500 ;
    LAYER M4 ;
      RECT 0.0000 230.2650 239.8000 239.6000 ;
      RECT 218.8850 230.1000 239.8000 230.2650 ;
      RECT 190.8300 230.1000 215.8850 230.2650 ;
      RECT 162.7750 230.1000 187.8300 230.2650 ;
      RECT 134.7200 230.1000 159.7750 230.2650 ;
      RECT 106.6650 230.1000 131.7200 230.2650 ;
      RECT 78.6100 230.1000 103.6650 230.2650 ;
      RECT 50.5550 230.1000 75.6100 230.2650 ;
      RECT 22.5000 230.1000 47.5550 230.2650 ;
      RECT 226.8850 9.5000 239.8000 230.1000 ;
      RECT 218.8850 9.5000 223.8850 230.1000 ;
      RECT 198.8300 9.5000 215.8850 230.1000 ;
      RECT 190.8300 9.5000 195.8300 230.1000 ;
      RECT 170.7750 9.5000 187.8300 230.1000 ;
      RECT 162.7750 9.5000 167.7750 230.1000 ;
      RECT 142.7200 9.5000 159.7750 230.1000 ;
      RECT 134.7200 9.5000 139.7200 230.1000 ;
      RECT 114.6650 9.5000 131.7200 230.1000 ;
      RECT 106.6650 9.5000 111.6650 230.1000 ;
      RECT 86.6100 9.5000 103.6650 230.1000 ;
      RECT 78.6100 9.5000 83.6100 230.1000 ;
      RECT 58.5550 9.5000 75.6100 230.1000 ;
      RECT 50.5550 9.5000 55.5550 230.1000 ;
      RECT 30.5000 9.5000 47.5550 230.1000 ;
      RECT 22.5000 9.5000 27.5000 230.1000 ;
      RECT 218.8850 9.3350 239.8000 9.5000 ;
      RECT 190.8300 9.3350 215.8850 9.5000 ;
      RECT 162.7750 9.3350 187.8300 9.5000 ;
      RECT 134.7200 9.3350 159.7750 9.5000 ;
      RECT 106.6650 9.3350 131.7200 9.5000 ;
      RECT 78.6100 9.3350 103.6650 9.5000 ;
      RECT 50.5550 9.3350 75.6100 9.5000 ;
      RECT 22.5000 9.3350 47.5550 9.5000 ;
      RECT 0.0000 9.3350 19.5000 230.2650 ;
      RECT 0.0000 0.0000 239.8000 9.3350 ;
  END
END sram_w16

END LIBRARY
