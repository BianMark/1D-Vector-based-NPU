##
## LEF for PtnCells ;
## created by Innovus v15.23-s045_1 on Fri Mar  7 16:13:28 2025
##

VERSION 5.8 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO fullchip
  CLASS BLOCK ;
  SIZE 554.0000 BY 551.0000 ;
  FOREIGN fullchip 0.0000 0.0000 ;
  ORIGIN 0 0 ;
  SYMMETRY X Y R90 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 275.7500 554.0000 275.8500 ;
    END
  END clk
  PIN mem_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 217.1500 0.5200 217.2500 ;
    END
  END mem_in[63]
  PIN mem_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 72.1500 0.5200 72.2500 ;
    END
  END mem_in[62]
  PIN mem_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 178.0500 0.0000 178.1500 0.5200 ;
    END
  END mem_in[61]
  PIN mem_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 117.9500 0.5200 118.0500 ;
    END
  END mem_in[60]
  PIN mem_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 215.9500 0.5200 216.0500 ;
    END
  END mem_in[59]
  PIN mem_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 205.1500 0.5200 205.2500 ;
    END
  END mem_in[58]
  PIN mem_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 86.1500 0.5200 86.2500 ;
    END
  END mem_in[57]
  PIN mem_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 186.5500 0.5200 186.6500 ;
    END
  END mem_in[56]
  PIN mem_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 91.5500 0.5200 91.6500 ;
    END
  END mem_in[55]
  PIN mem_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 134.1500 0.5200 134.2500 ;
    END
  END mem_in[54]
  PIN mem_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 100.6500 0.0000 100.7500 0.5200 ;
    END
  END mem_in[53]
  PIN mem_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.8500 0.0000 164.9500 0.5200 ;
    END
  END mem_in[52]
  PIN mem_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 185.2500 0.0000 185.3500 0.5200 ;
    END
  END mem_in[51]
  PIN mem_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 194.2500 0.0000 194.3500 0.5200 ;
    END
  END mem_in[50]
  PIN mem_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 106.4500 0.0000 106.5500 0.5200 ;
    END
  END mem_in[49]
  PIN mem_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 123.0500 0.0000 123.1500 0.5200 ;
    END
  END mem_in[48]
  PIN mem_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 201.1500 0.5200 201.2500 ;
    END
  END mem_in[47]
  PIN mem_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 216.5500 0.5200 216.6500 ;
    END
  END mem_in[46]
  PIN mem_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 192.4500 0.0000 192.5500 0.5200 ;
    END
  END mem_in[45]
  PIN mem_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 215.5500 0.5200 215.6500 ;
    END
  END mem_in[44]
  PIN mem_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 209.7500 0.5200 209.8500 ;
    END
  END mem_in[43]
  PIN mem_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 194.9500 0.5200 195.0500 ;
    END
  END mem_in[42]
  PIN mem_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 75.6500 0.0000 75.7500 0.5200 ;
    END
  END mem_in[41]
  PIN mem_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 119.6500 0.0000 119.7500 0.5200 ;
    END
  END mem_in[40]
  PIN mem_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 211.1500 0.5200 211.2500 ;
    END
  END mem_in[39]
  PIN mem_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 134.0500 0.0000 134.1500 0.5200 ;
    END
  END mem_in[38]
  PIN mem_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 105.8500 0.0000 105.9500 0.5200 ;
    END
  END mem_in[37]
  PIN mem_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 205.7500 0.5200 205.8500 ;
    END
  END mem_in[36]
  PIN mem_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 96.1500 0.5200 96.2500 ;
    END
  END mem_in[35]
  PIN mem_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 127.6500 0.0000 127.7500 0.5200 ;
    END
  END mem_in[34]
  PIN mem_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 210.1500 0.5200 210.2500 ;
    END
  END mem_in[33]
  PIN mem_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 104.2500 0.0000 104.3500 0.5200 ;
    END
  END mem_in[32]
  PIN mem_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 187.4500 0.0000 187.5500 0.5200 ;
    END
  END mem_in[31]
  PIN mem_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 191.8500 0.0000 191.9500 0.5200 ;
    END
  END mem_in[30]
  PIN mem_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 197.9500 0.5200 198.0500 ;
    END
  END mem_in[29]
  PIN mem_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 131.3500 0.5200 131.4500 ;
    END
  END mem_in[28]
  PIN mem_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 181.6500 0.0000 181.7500 0.5200 ;
    END
  END mem_in[27]
  PIN mem_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 167.8500 0.0000 167.9500 0.5200 ;
    END
  END mem_in[26]
  PIN mem_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 219.3500 0.5200 219.4500 ;
    END
  END mem_in[25]
  PIN mem_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 210.5500 0.5200 210.6500 ;
    END
  END mem_in[24]
  PIN mem_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 209.3500 0.5200 209.4500 ;
    END
  END mem_in[23]
  PIN mem_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 65.4500 0.0000 65.5500 0.5200 ;
    END
  END mem_in[22]
  PIN mem_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 91.9500 0.5200 92.0500 ;
    END
  END mem_in[21]
  PIN mem_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 71.7500 0.5200 71.8500 ;
    END
  END mem_in[20]
  PIN mem_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 191.5500 0.5200 191.6500 ;
    END
  END mem_in[19]
  PIN mem_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 227.7500 0.5200 227.8500 ;
    END
  END mem_in[18]
  PIN mem_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 169.2500 0.0000 169.3500 0.5200 ;
    END
  END mem_in[17]
  PIN mem_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 213.1500 0.5200 213.2500 ;
    END
  END mem_in[16]
  PIN mem_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 73.7500 0.5200 73.8500 ;
    END
  END mem_in[15]
  PIN mem_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 220.3500 0.5200 220.4500 ;
    END
  END mem_in[14]
  PIN mem_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 57.1500 0.5200 57.2500 ;
    END
  END mem_in[13]
  PIN mem_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 171.2500 0.0000 171.3500 0.5200 ;
    END
  END mem_in[12]
  PIN mem_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 204.1500 0.5200 204.2500 ;
    END
  END mem_in[11]
  PIN mem_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 164.2500 0.0000 164.3500 0.5200 ;
    END
  END mem_in[10]
  PIN mem_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 133.0500 0.0000 133.1500 0.5200 ;
    END
  END mem_in[9]
  PIN mem_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 77.6500 0.0000 77.7500 0.5200 ;
    END
  END mem_in[8]
  PIN mem_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 203.3500 0.5200 203.4500 ;
    END
  END mem_in[7]
  PIN mem_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 76.1500 0.5200 76.2500 ;
    END
  END mem_in[6]
  PIN mem_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 72.7500 0.5200 72.8500 ;
    END
  END mem_in[5]
  PIN mem_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 164.8500 0.0000 164.9500 0.5200 ;
    END
  END mem_in[4]
  PIN mem_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 208.3500 0.5200 208.4500 ;
    END
  END mem_in[3]
  PIN mem_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 193.5500 0.5200 193.6500 ;
    END
  END mem_in[2]
  PIN mem_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 215.1500 0.5200 215.2500 ;
    END
  END mem_in[1]
  PIN mem_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 71.3500 0.5200 71.4500 ;
    END
  END mem_in[0]
  PIN inst[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 304.7500 554.0000 304.8500 ;
    END
  END inst[16]
  PIN inst[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 198.3500 0.5200 198.4500 ;
    END
  END inst[15]
  PIN inst[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 195.9500 0.5200 196.0500 ;
    END
  END inst[14]
  PIN inst[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 195.3500 0.5200 195.4500 ;
    END
  END inst[13]
  PIN inst[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 198.7500 0.5200 198.8500 ;
    END
  END inst[12]
  PIN inst[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 268.2500 550.4800 268.3500 551.0000 ;
    END
  END inst[11]
  PIN inst[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 269.2500 550.4800 269.3500 551.0000 ;
    END
  END inst[10]
  PIN inst[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.2500 550.4800 280.3500 551.0000 ;
    END
  END inst[9]
  PIN inst[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 280.8500 550.4800 280.9500 551.0000 ;
    END
  END inst[8]
  PIN inst[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 282.4500 0.0000 282.5500 0.5200 ;
    END
  END inst[7]
  PIN inst[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 120.3500 0.5200 120.4500 ;
    END
  END inst[6]
  PIN inst[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 523.7500 0.5200 523.8500 ;
    END
  END inst[5]
  PIN inst[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 523.3500 0.5200 523.4500 ;
    END
  END inst[4]
  PIN inst[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 12.4500 550.4800 12.5500 551.0000 ;
    END
  END inst[3]
  PIN inst[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 13.2500 550.4800 13.3500 551.0000 ;
    END
  END inst[2]
  PIN inst[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 530.9500 0.5200 531.0500 ;
    END
  END inst[1]
  PIN inst[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 0.0000 531.9500 0.5200 532.0500 ;
    END
  END inst[0]
  PIN reset
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 276.6500 550.4800 276.7500 551.0000 ;
    END
  END reset
  PIN out[159]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 344.1500 554.0000 344.2500 ;
    END
  END out[159]
  PIN out[158]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 338.1500 554.0000 338.2500 ;
    END
  END out[158]
  PIN out[157]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 374.1500 554.0000 374.2500 ;
    END
  END out[157]
  PIN out[156]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 370.5500 554.0000 370.6500 ;
    END
  END out[156]
  PIN out[155]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 329.7500 554.0000 329.8500 ;
    END
  END out[155]
  PIN out[154]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 308.1500 554.0000 308.2500 ;
    END
  END out[154]
  PIN out[153]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 334.5500 554.0000 334.6500 ;
    END
  END out[153]
  PIN out[152]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 399.3500 554.0000 399.4500 ;
    END
  END out[152]
  PIN out[151]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 383.7500 554.0000 383.8500 ;
    END
  END out[151]
  PIN out[150]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 333.3500 554.0000 333.4500 ;
    END
  END out[150]
  PIN out[149]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 417.3500 554.0000 417.4500 ;
    END
  END out[149]
  PIN out[148]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 348.9500 554.0000 349.0500 ;
    END
  END out[148]
  PIN out[147]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 423.3500 554.0000 423.4500 ;
    END
  END out[147]
  PIN out[146]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 329.3500 554.0000 329.4500 ;
    END
  END out[146]
  PIN out[145]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 269.7500 554.0000 269.8500 ;
    END
  END out[145]
  PIN out[144]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 359.7500 554.0000 359.8500 ;
    END
  END out[144]
  PIN out[143]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 307.7500 554.0000 307.8500 ;
    END
  END out[143]
  PIN out[142]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 293.7500 554.0000 293.8500 ;
    END
  END out[142]
  PIN out[141]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 420.9500 554.0000 421.0500 ;
    END
  END out[141]
  PIN out[140]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 345.3500 554.0000 345.4500 ;
    END
  END out[140]
  PIN out[139]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 394.5500 554.0000 394.6500 ;
    END
  END out[139]
  PIN out[138]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 456.9500 554.0000 457.0500 ;
    END
  END out[138]
  PIN out[137]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 402.9500 554.0000 403.0500 ;
    END
  END out[137]
  PIN out[136]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 473.7500 554.0000 473.8500 ;
    END
  END out[136]
  PIN out[135]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 498.9500 554.0000 499.0500 ;
    END
  END out[135]
  PIN out[134]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 480.9500 554.0000 481.0500 ;
    END
  END out[134]
  PIN out[133]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 419.7500 554.0000 419.8500 ;
    END
  END out[133]
  PIN out[132]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 373.7500 554.0000 373.8500 ;
    END
  END out[132]
  PIN out[131]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 464.1500 554.0000 464.2500 ;
    END
  END out[131]
  PIN out[130]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 460.4500 550.4800 460.5500 551.0000 ;
    END
  END out[130]
  PIN out[129]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 416.1500 554.0000 416.2500 ;
    END
  END out[129]
  PIN out[128]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 532.5500 554.0000 532.6500 ;
    END
  END out[128]
  PIN out[127]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 420.5500 554.0000 420.6500 ;
    END
  END out[127]
  PIN out[126]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 510.6500 550.4800 510.7500 551.0000 ;
    END
  END out[126]
  PIN out[125]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 524.1500 554.0000 524.2500 ;
    END
  END out[125]
  PIN out[124]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 437.7500 554.0000 437.8500 ;
    END
  END out[124]
  PIN out[123]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 438.9500 554.0000 439.0500 ;
    END
  END out[123]
  PIN out[122]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 495.3500 554.0000 495.4500 ;
    END
  END out[122]
  PIN out[121]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 442.5500 554.0000 442.6500 ;
    END
  END out[121]
  PIN out[120]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 380.1500 554.0000 380.2500 ;
    END
  END out[120]
  PIN out[119]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 264.9500 554.0000 265.0500 ;
    END
  END out[119]
  PIN out[118]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 192.9500 554.0000 193.0500 ;
    END
  END out[118]
  PIN out[117]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 272.1500 554.0000 272.2500 ;
    END
  END out[117]
  PIN out[116]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 219.3500 554.0000 219.4500 ;
    END
  END out[116]
  PIN out[115]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 268.5500 554.0000 268.6500 ;
    END
  END out[115]
  PIN out[114]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 261.3500 554.0000 261.4500 ;
    END
  END out[114]
  PIN out[113]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 293.3500 554.0000 293.4500 ;
    END
  END out[113]
  PIN out[112]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 192.5500 554.0000 192.6500 ;
    END
  END out[112]
  PIN out[111]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 280.5500 554.0000 280.6500 ;
    END
  END out[111]
  PIN out[110]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 322.5500 554.0000 322.6500 ;
    END
  END out[110]
  PIN out[109]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 128.1500 554.0000 128.2500 ;
    END
  END out[109]
  PIN out[108]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 232.5500 554.0000 232.6500 ;
    END
  END out[108]
  PIN out[107]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 215.7500 554.0000 215.8500 ;
    END
  END out[107]
  PIN out[106]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 341.7500 554.0000 341.8500 ;
    END
  END out[106]
  PIN out[105]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 271.7500 554.0000 271.8500 ;
    END
  END out[105]
  PIN out[104]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 185.7500 554.0000 185.8500 ;
    END
  END out[104]
  PIN out[103]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 251.7500 554.0000 251.8500 ;
    END
  END out[103]
  PIN out[102]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 266.1500 554.0000 266.2500 ;
    END
  END out[102]
  PIN out[101]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 282.9500 554.0000 283.0500 ;
    END
  END out[101]
  PIN out[100]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 260.9500 554.0000 261.0500 ;
    END
  END out[100]
  PIN out[99]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 519.0500 550.4800 519.1500 551.0000 ;
    END
  END out[99]
  PIN out[98]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 498.5500 554.0000 498.6500 ;
    END
  END out[98]
  PIN out[97]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 500.1500 554.0000 500.2500 ;
    END
  END out[97]
  PIN out[96]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 536.1500 554.0000 536.2500 ;
    END
  END out[96]
  PIN out[95]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 477.2500 550.4800 477.3500 551.0000 ;
    END
  END out[95]
  PIN out[94]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 443.6500 550.4800 443.7500 551.0000 ;
    END
  END out[94]
  PIN out[93]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 513.3500 554.0000 513.4500 ;
    END
  END out[93]
  PIN out[92]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 538.5500 554.0000 538.6500 ;
    END
  END out[92]
  PIN out[91]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 455.7500 554.0000 455.8500 ;
    END
  END out[91]
  PIN out[90]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 531.3500 554.0000 531.4500 ;
    END
  END out[90]
  PIN out[89]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 534.9500 554.0000 535.0500 ;
    END
  END out[89]
  PIN out[88]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 528.9500 554.0000 529.0500 ;
    END
  END out[88]
  PIN out[87]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 492.9500 554.0000 493.0500 ;
    END
  END out[87]
  PIN out[86]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 462.9500 554.0000 463.0500 ;
    END
  END out[86]
  PIN out[85]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 530.9500 554.0000 531.0500 ;
    END
  END out[85]
  PIN out[84]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 459.3500 554.0000 459.4500 ;
    END
  END out[84]
  PIN out[83]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 496.5500 554.0000 496.6500 ;
    END
  END out[83]
  PIN out[82]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 426.9500 554.0000 427.0500 ;
    END
  END out[82]
  PIN out[81]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 484.5500 554.0000 484.6500 ;
    END
  END out[81]
  PIN out[80]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 512.9500 554.0000 513.0500 ;
    END
  END out[80]
  PIN out[79]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 351.3500 554.0000 351.4500 ;
    END
  END out[79]
  PIN out[78]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 499.3500 554.0000 499.4500 ;
    END
  END out[78]
  PIN out[77]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 444.9500 554.0000 445.0500 ;
    END
  END out[77]
  PIN out[76]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 502.2500 550.4800 502.3500 551.0000 ;
    END
  END out[76]
  PIN out[75]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 428.1500 554.0000 428.2500 ;
    END
  END out[75]
  PIN out[74]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 424.5500 554.0000 424.6500 ;
    END
  END out[74]
  PIN out[73]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 398.1500 554.0000 398.2500 ;
    END
  END out[73]
  PIN out[72]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 225.3500 554.0000 225.4500 ;
    END
  END out[72]
  PIN out[71]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 416.9500 554.0000 417.0500 ;
    END
  END out[71]
  PIN out[70]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 521.7500 554.0000 521.8500 ;
    END
  END out[70]
  PIN out[69]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 401.7500 554.0000 401.8500 ;
    END
  END out[69]
  PIN out[68]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 503.7500 554.0000 503.8500 ;
    END
  END out[68]
  PIN out[67]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 519.0500 550.4800 519.1500 551.0000 ;
    END
  END out[67]
  PIN out[66]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 377.7500 554.0000 377.8500 ;
    END
  END out[66]
  PIN out[65]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 532.1500 554.0000 532.2500 ;
    END
  END out[65]
  PIN out[64]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 427.7500 554.0000 427.8500 ;
    END
  END out[64]
  PIN out[63]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 395.7500 554.0000 395.8500 ;
    END
  END out[63]
  PIN out[62]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 460.5500 554.0000 460.6500 ;
    END
  END out[62]
  PIN out[61]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 352.5500 554.0000 352.6500 ;
    END
  END out[61]
  PIN out[60]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 502.5500 554.0000 502.6500 ;
    END
  END out[60]
  PIN out[59]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 492.5500 554.0000 492.6500 ;
    END
  END out[59]
  PIN out[58]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 527.4500 550.4800 527.5500 551.0000 ;
    END
  END out[58]
  PIN out[57]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 473.3500 554.0000 473.4500 ;
    END
  END out[57]
  PIN out[56]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 535.8500 550.4800 535.9500 551.0000 ;
    END
  END out[56]
  PIN out[55]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 535.8500 550.4800 535.9500 551.0000 ;
    END
  END out[55]
  PIN out[54]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 447.6500 550.4800 447.7500 551.0000 ;
    END
  END out[54]
  PIN out[53]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 467.7500 554.0000 467.8500 ;
    END
  END out[53]
  PIN out[52]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 527.7500 554.0000 527.8500 ;
    END
  END out[52]
  PIN out[51]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 539.7500 554.0000 539.8500 ;
    END
  END out[51]
  PIN out[50]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 419.3500 554.0000 419.4500 ;
    END
  END out[50]
  PIN out[49]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 510.6500 550.4800 510.7500 551.0000 ;
    END
  END out[49]
  PIN out[48]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 525.3500 554.0000 525.4500 ;
    END
  END out[48]
  PIN out[47]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 482.1500 554.0000 482.2500 ;
    END
  END out[47]
  PIN out[46]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 474.1500 554.0000 474.2500 ;
    END
  END out[46]
  PIN out[45]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 510.2500 550.4800 510.3500 551.0000 ;
    END
  END out[45]
  PIN out[44]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 511.0500 550.4800 511.1500 551.0000 ;
    END
  END out[44]
  PIN out[43]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 458.9500 554.0000 459.0500 ;
    END
  END out[43]
  PIN out[42]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 438.5500 554.0000 438.6500 ;
    END
  END out[42]
  PIN out[41]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 524.9500 554.0000 525.0500 ;
    END
  END out[41]
  PIN out[40]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 498.1500 554.0000 498.2500 ;
    END
  END out[40]
  PIN out[39]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 218.9500 554.0000 219.0500 ;
    END
  END out[39]
  PIN out[38]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 107.7500 554.0000 107.8500 ;
    END
  END out[38]
  PIN out[37]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 219.7500 554.0000 219.8500 ;
    END
  END out[37]
  PIN out[36]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 250.5500 554.0000 250.6500 ;
    END
  END out[36]
  PIN out[35]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 257.7500 554.0000 257.8500 ;
    END
  END out[35]
  PIN out[34]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 294.9500 554.0000 295.0500 ;
    END
  END out[34]
  PIN out[33]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 273.3500 554.0000 273.4500 ;
    END
  END out[33]
  PIN out[32]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 243.3500 554.0000 243.4500 ;
    END
  END out[32]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 194.1500 554.0000 194.2500 ;
    END
  END out[31]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 272.9500 554.0000 273.0500 ;
    END
  END out[30]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 240.9500 554.0000 241.0500 ;
    END
  END out[29]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 255.3500 554.0000 255.4500 ;
    END
  END out[28]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 248.1500 554.0000 248.2500 ;
    END
  END out[27]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 218.1500 554.0000 218.2500 ;
    END
  END out[26]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 215.3500 554.0000 215.4500 ;
    END
  END out[25]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 250.1500 554.0000 250.2500 ;
    END
  END out[24]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 217.7500 554.0000 217.8500 ;
    END
  END out[23]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 239.7500 554.0000 239.8500 ;
    END
  END out[22]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 237.3500 554.0000 237.4500 ;
    END
  END out[21]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 172.5500 554.0000 172.6500 ;
    END
  END out[20]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 224.9500 554.0000 225.0500 ;
    END
  END out[19]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 485.6500 0.0000 485.7500 0.5200 ;
    END
  END out[18]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 435.2500 0.0000 435.3500 0.5200 ;
    END
  END out[17]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 485.6500 0.0000 485.7500 0.5200 ;
    END
  END out[16]
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 340.5500 554.0000 340.6500 ;
    END
  END out[15]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 302.1500 554.0000 302.2500 ;
    END
  END out[14]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 140.1500 554.0000 140.2500 ;
    END
  END out[13]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 294.1500 554.0000 294.2500 ;
    END
  END out[12]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 410.4500 0.0000 410.5500 0.5200 ;
    END
  END out[11]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 261.7500 554.0000 261.8500 ;
    END
  END out[10]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 347.7500 554.0000 347.8500 ;
    END
  END out[9]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 427.0500 0.0000 427.1500 0.5200 ;
    END
  END out[8]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 146.1500 554.0000 146.2500 ;
    END
  END out[7]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M2 ;
        RECT 477.2500 0.0000 477.3500 0.5200 ;
    END
  END out[6]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 222.9500 554.0000 223.0500 ;
    END
  END out[5]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 240.5500 554.0000 240.6500 ;
    END
  END out[4]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 336.9500 554.0000 337.0500 ;
    END
  END out[3]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 347.3500 554.0000 347.4500 ;
    END
  END out[2]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M4 ;
        RECT 477.2500 0.0000 477.3500 0.5200 ;
    END
  END out[1]
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER M3 ;
        RECT 553.4800 113.7500 554.0000 113.8500 ;
    END
  END out[0]
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 196.3300 6.0000 198.3300 545.0000 ;
        RECT 168.2750 6.0000 170.2750 545.0000 ;
        RECT 140.2200 6.0000 142.2200 545.0000 ;
        RECT 112.1650 6.0000 114.1650 545.0000 ;
        RECT 84.1100 6.0000 86.1100 545.0000 ;
        RECT 56.0550 6.0000 58.0550 545.0000 ;
        RECT 28.0000 6.0000 30.0000 545.0000 ;
        RECT 224.3850 6.0000 226.3850 545.0000 ;
        RECT 252.4400 6.0000 254.4400 545.0000 ;
        RECT 280.4950 6.0000 282.4950 545.0000 ;
        RECT 308.5500 6.0000 310.5500 545.0000 ;
        RECT 336.6050 6.0000 338.6050 545.0000 ;
        RECT 364.6600 6.0000 366.6600 545.0000 ;
        RECT 392.7150 6.0000 394.7150 545.0000 ;
        RECT 420.7700 6.0000 422.7700 545.0000 ;
        RECT 448.8250 6.0000 450.8250 545.0000 ;
        RECT 476.8800 6.0000 478.8800 545.0000 ;
        RECT 504.9350 6.0000 506.9350 545.0000 ;
        RECT 532.9900 6.0000 534.9900 545.0000 ;
    END
# end of P/G power stripe data as pin

  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;

# P/G power stripe data as pin
    PORT
      LAYER M4 ;
        RECT 272.4950 1.0000 274.4950 550.0000 ;
        RECT 244.4400 1.0000 246.4400 550.0000 ;
        RECT 216.3850 1.0000 218.3850 550.0000 ;
        RECT 188.3300 1.0000 190.3300 550.0000 ;
        RECT 160.2750 1.0000 162.2750 550.0000 ;
        RECT 132.2200 1.0000 134.2200 550.0000 ;
        RECT 104.1650 1.0000 106.1650 550.0000 ;
        RECT 76.1100 1.0000 78.1100 550.0000 ;
        RECT 48.0550 1.0000 50.0550 550.0000 ;
        RECT 20.0000 1.0000 22.0000 550.0000 ;
        RECT 524.9900 1.0000 526.9900 550.0000 ;
        RECT 496.9350 1.0000 498.9350 550.0000 ;
        RECT 468.8800 1.0000 470.8800 550.0000 ;
        RECT 440.8250 1.0000 442.8250 550.0000 ;
        RECT 412.7700 1.0000 414.7700 550.0000 ;
        RECT 384.7150 1.0000 386.7150 550.0000 ;
        RECT 356.6600 1.0000 358.6600 550.0000 ;
        RECT 328.6050 1.0000 330.6050 550.0000 ;
        RECT 300.5500 1.0000 302.5500 550.0000 ;
    END
# end of P/G power stripe data as pin

  END VDD
  OBS
    LAYER M1 ;
      RECT 0.0000 0.0000 554.0000 551.0000 ;
    LAYER M2 ;
      RECT 536.0500 550.3800 554.0000 551.0000 ;
      RECT 527.6500 550.3800 535.7500 551.0000 ;
      RECT 519.2500 550.3800 527.3500 551.0000 ;
      RECT 511.2500 550.3800 518.9500 551.0000 ;
      RECT 510.8500 550.3800 510.9500 551.0000 ;
      RECT 510.4500 550.3800 510.5500 551.0000 ;
      RECT 502.4500 550.3800 510.1500 551.0000 ;
      RECT 477.4500 550.3800 502.1500 551.0000 ;
      RECT 460.6500 550.3800 477.1500 551.0000 ;
      RECT 447.8500 550.3800 460.3500 551.0000 ;
      RECT 443.8500 550.3800 447.5500 551.0000 ;
      RECT 281.0500 550.3800 443.5500 551.0000 ;
      RECT 280.4500 550.3800 280.7500 551.0000 ;
      RECT 276.8500 550.3800 280.1500 551.0000 ;
      RECT 269.4500 550.3800 276.5500 551.0000 ;
      RECT 268.4500 550.3800 269.1500 551.0000 ;
      RECT 13.4500 550.3800 268.1500 551.0000 ;
      RECT 12.6500 550.3800 13.1500 551.0000 ;
      RECT 0.0000 550.3800 12.3500 551.0000 ;
      RECT 0.0000 0.6200 554.0000 550.3800 ;
      RECT 485.8500 0.0000 554.0000 0.6200 ;
      RECT 477.4500 0.0000 485.5500 0.6200 ;
      RECT 435.4500 0.0000 477.1500 0.6200 ;
      RECT 427.2500 0.0000 435.1500 0.6200 ;
      RECT 410.6500 0.0000 426.9500 0.6200 ;
      RECT 282.6500 0.0000 410.3500 0.6200 ;
      RECT 194.4500 0.0000 282.3500 0.6200 ;
      RECT 192.6500 0.0000 194.1500 0.6200 ;
      RECT 192.0500 0.0000 192.3500 0.6200 ;
      RECT 187.6500 0.0000 191.7500 0.6200 ;
      RECT 185.4500 0.0000 187.3500 0.6200 ;
      RECT 181.8500 0.0000 185.1500 0.6200 ;
      RECT 178.2500 0.0000 181.5500 0.6200 ;
      RECT 171.4500 0.0000 177.9500 0.6200 ;
      RECT 169.4500 0.0000 171.1500 0.6200 ;
      RECT 168.0500 0.0000 169.1500 0.6200 ;
      RECT 165.0500 0.0000 167.7500 0.6200 ;
      RECT 164.4500 0.0000 164.7500 0.6200 ;
      RECT 134.2500 0.0000 164.1500 0.6200 ;
      RECT 133.2500 0.0000 133.9500 0.6200 ;
      RECT 127.8500 0.0000 132.9500 0.6200 ;
      RECT 123.2500 0.0000 127.5500 0.6200 ;
      RECT 119.8500 0.0000 122.9500 0.6200 ;
      RECT 106.6500 0.0000 119.5500 0.6200 ;
      RECT 106.0500 0.0000 106.3500 0.6200 ;
      RECT 104.4500 0.0000 105.7500 0.6200 ;
      RECT 100.8500 0.0000 104.1500 0.6200 ;
      RECT 77.8500 0.0000 100.5500 0.6200 ;
      RECT 75.8500 0.0000 77.5500 0.6200 ;
      RECT 65.6500 0.0000 75.5500 0.6200 ;
      RECT 0.0000 0.0000 65.3500 0.6200 ;
    LAYER M3 ;
      RECT 0.0000 539.9500 554.0000 551.0000 ;
      RECT 0.0000 539.6500 553.3800 539.9500 ;
      RECT 0.0000 538.7500 554.0000 539.6500 ;
      RECT 0.0000 538.4500 553.3800 538.7500 ;
      RECT 0.0000 536.3500 554.0000 538.4500 ;
      RECT 0.0000 536.0500 553.3800 536.3500 ;
      RECT 0.0000 535.1500 554.0000 536.0500 ;
      RECT 0.0000 534.8500 553.3800 535.1500 ;
      RECT 0.0000 532.7500 554.0000 534.8500 ;
      RECT 0.0000 532.4500 553.3800 532.7500 ;
      RECT 0.0000 532.3500 554.0000 532.4500 ;
      RECT 0.0000 532.1500 553.3800 532.3500 ;
      RECT 0.6200 532.0500 553.3800 532.1500 ;
      RECT 0.6200 531.8500 554.0000 532.0500 ;
      RECT 0.0000 531.5500 554.0000 531.8500 ;
      RECT 0.0000 531.2500 553.3800 531.5500 ;
      RECT 0.0000 531.1500 554.0000 531.2500 ;
      RECT 0.6200 530.8500 553.3800 531.1500 ;
      RECT 0.0000 529.1500 554.0000 530.8500 ;
      RECT 0.0000 528.8500 553.3800 529.1500 ;
      RECT 0.0000 527.9500 554.0000 528.8500 ;
      RECT 0.0000 527.6500 553.3800 527.9500 ;
      RECT 0.0000 525.5500 554.0000 527.6500 ;
      RECT 0.0000 525.2500 553.3800 525.5500 ;
      RECT 0.0000 525.1500 554.0000 525.2500 ;
      RECT 0.0000 524.8500 553.3800 525.1500 ;
      RECT 0.0000 524.3500 554.0000 524.8500 ;
      RECT 0.0000 524.0500 553.3800 524.3500 ;
      RECT 0.0000 523.9500 554.0000 524.0500 ;
      RECT 0.6200 523.6500 554.0000 523.9500 ;
      RECT 0.0000 523.5500 554.0000 523.6500 ;
      RECT 0.6200 523.2500 554.0000 523.5500 ;
      RECT 0.0000 521.9500 554.0000 523.2500 ;
      RECT 0.0000 521.6500 553.3800 521.9500 ;
      RECT 0.0000 513.5500 554.0000 521.6500 ;
      RECT 0.0000 513.2500 553.3800 513.5500 ;
      RECT 0.0000 513.1500 554.0000 513.2500 ;
      RECT 0.0000 512.8500 553.3800 513.1500 ;
      RECT 0.0000 503.9500 554.0000 512.8500 ;
      RECT 0.0000 503.6500 553.3800 503.9500 ;
      RECT 0.0000 502.7500 554.0000 503.6500 ;
      RECT 0.0000 502.4500 553.3800 502.7500 ;
      RECT 0.0000 500.3500 554.0000 502.4500 ;
      RECT 0.0000 500.0500 553.3800 500.3500 ;
      RECT 0.0000 499.5500 554.0000 500.0500 ;
      RECT 0.0000 499.2500 553.3800 499.5500 ;
      RECT 0.0000 499.1500 554.0000 499.2500 ;
      RECT 0.0000 498.8500 553.3800 499.1500 ;
      RECT 0.0000 498.7500 554.0000 498.8500 ;
      RECT 0.0000 498.4500 553.3800 498.7500 ;
      RECT 0.0000 498.3500 554.0000 498.4500 ;
      RECT 0.0000 498.0500 553.3800 498.3500 ;
      RECT 0.0000 496.7500 554.0000 498.0500 ;
      RECT 0.0000 496.4500 553.3800 496.7500 ;
      RECT 0.0000 495.5500 554.0000 496.4500 ;
      RECT 0.0000 495.2500 553.3800 495.5500 ;
      RECT 0.0000 493.1500 554.0000 495.2500 ;
      RECT 0.0000 492.8500 553.3800 493.1500 ;
      RECT 0.0000 492.7500 554.0000 492.8500 ;
      RECT 0.0000 492.4500 553.3800 492.7500 ;
      RECT 0.0000 484.7500 554.0000 492.4500 ;
      RECT 0.0000 484.4500 553.3800 484.7500 ;
      RECT 0.0000 482.3500 554.0000 484.4500 ;
      RECT 0.0000 482.0500 553.3800 482.3500 ;
      RECT 0.0000 481.1500 554.0000 482.0500 ;
      RECT 0.0000 480.8500 553.3800 481.1500 ;
      RECT 0.0000 474.3500 554.0000 480.8500 ;
      RECT 0.0000 474.0500 553.3800 474.3500 ;
      RECT 0.0000 473.9500 554.0000 474.0500 ;
      RECT 0.0000 473.6500 553.3800 473.9500 ;
      RECT 0.0000 473.5500 554.0000 473.6500 ;
      RECT 0.0000 473.2500 553.3800 473.5500 ;
      RECT 0.0000 467.9500 554.0000 473.2500 ;
      RECT 0.0000 467.6500 553.3800 467.9500 ;
      RECT 0.0000 464.3500 554.0000 467.6500 ;
      RECT 0.0000 464.0500 553.3800 464.3500 ;
      RECT 0.0000 463.1500 554.0000 464.0500 ;
      RECT 0.0000 462.8500 553.3800 463.1500 ;
      RECT 0.0000 460.7500 554.0000 462.8500 ;
      RECT 0.0000 460.4500 553.3800 460.7500 ;
      RECT 0.0000 459.5500 554.0000 460.4500 ;
      RECT 0.0000 459.2500 553.3800 459.5500 ;
      RECT 0.0000 459.1500 554.0000 459.2500 ;
      RECT 0.0000 458.8500 553.3800 459.1500 ;
      RECT 0.0000 457.1500 554.0000 458.8500 ;
      RECT 0.0000 456.8500 553.3800 457.1500 ;
      RECT 0.0000 455.9500 554.0000 456.8500 ;
      RECT 0.0000 455.6500 553.3800 455.9500 ;
      RECT 0.0000 445.1500 554.0000 455.6500 ;
      RECT 0.0000 444.8500 553.3800 445.1500 ;
      RECT 0.0000 442.7500 554.0000 444.8500 ;
      RECT 0.0000 442.4500 553.3800 442.7500 ;
      RECT 0.0000 439.1500 554.0000 442.4500 ;
      RECT 0.0000 438.8500 553.3800 439.1500 ;
      RECT 0.0000 438.7500 554.0000 438.8500 ;
      RECT 0.0000 438.4500 553.3800 438.7500 ;
      RECT 0.0000 437.9500 554.0000 438.4500 ;
      RECT 0.0000 437.6500 553.3800 437.9500 ;
      RECT 0.0000 428.3500 554.0000 437.6500 ;
      RECT 0.0000 428.0500 553.3800 428.3500 ;
      RECT 0.0000 427.9500 554.0000 428.0500 ;
      RECT 0.0000 427.6500 553.3800 427.9500 ;
      RECT 0.0000 427.1500 554.0000 427.6500 ;
      RECT 0.0000 426.8500 553.3800 427.1500 ;
      RECT 0.0000 424.7500 554.0000 426.8500 ;
      RECT 0.0000 424.4500 553.3800 424.7500 ;
      RECT 0.0000 423.5500 554.0000 424.4500 ;
      RECT 0.0000 423.2500 553.3800 423.5500 ;
      RECT 0.0000 421.1500 554.0000 423.2500 ;
      RECT 0.0000 420.8500 553.3800 421.1500 ;
      RECT 0.0000 420.7500 554.0000 420.8500 ;
      RECT 0.0000 420.4500 553.3800 420.7500 ;
      RECT 0.0000 419.9500 554.0000 420.4500 ;
      RECT 0.0000 419.6500 553.3800 419.9500 ;
      RECT 0.0000 419.5500 554.0000 419.6500 ;
      RECT 0.0000 419.2500 553.3800 419.5500 ;
      RECT 0.0000 417.5500 554.0000 419.2500 ;
      RECT 0.0000 417.2500 553.3800 417.5500 ;
      RECT 0.0000 417.1500 554.0000 417.2500 ;
      RECT 0.0000 416.8500 553.3800 417.1500 ;
      RECT 0.0000 416.3500 554.0000 416.8500 ;
      RECT 0.0000 416.0500 553.3800 416.3500 ;
      RECT 0.0000 403.1500 554.0000 416.0500 ;
      RECT 0.0000 402.8500 553.3800 403.1500 ;
      RECT 0.0000 401.9500 554.0000 402.8500 ;
      RECT 0.0000 401.6500 553.3800 401.9500 ;
      RECT 0.0000 399.5500 554.0000 401.6500 ;
      RECT 0.0000 399.2500 553.3800 399.5500 ;
      RECT 0.0000 398.3500 554.0000 399.2500 ;
      RECT 0.0000 398.0500 553.3800 398.3500 ;
      RECT 0.0000 395.9500 554.0000 398.0500 ;
      RECT 0.0000 395.6500 553.3800 395.9500 ;
      RECT 0.0000 394.7500 554.0000 395.6500 ;
      RECT 0.0000 394.4500 553.3800 394.7500 ;
      RECT 0.0000 383.9500 554.0000 394.4500 ;
      RECT 0.0000 383.6500 553.3800 383.9500 ;
      RECT 0.0000 380.3500 554.0000 383.6500 ;
      RECT 0.0000 380.0500 553.3800 380.3500 ;
      RECT 0.0000 377.9500 554.0000 380.0500 ;
      RECT 0.0000 377.6500 553.3800 377.9500 ;
      RECT 0.0000 374.3500 554.0000 377.6500 ;
      RECT 0.0000 374.0500 553.3800 374.3500 ;
      RECT 0.0000 373.9500 554.0000 374.0500 ;
      RECT 0.0000 373.6500 553.3800 373.9500 ;
      RECT 0.0000 370.7500 554.0000 373.6500 ;
      RECT 0.0000 370.4500 553.3800 370.7500 ;
      RECT 0.0000 359.9500 554.0000 370.4500 ;
      RECT 0.0000 359.6500 553.3800 359.9500 ;
      RECT 0.0000 352.7500 554.0000 359.6500 ;
      RECT 0.0000 352.4500 553.3800 352.7500 ;
      RECT 0.0000 351.5500 554.0000 352.4500 ;
      RECT 0.0000 351.2500 553.3800 351.5500 ;
      RECT 0.0000 349.1500 554.0000 351.2500 ;
      RECT 0.0000 348.8500 553.3800 349.1500 ;
      RECT 0.0000 347.9500 554.0000 348.8500 ;
      RECT 0.0000 347.6500 553.3800 347.9500 ;
      RECT 0.0000 347.5500 554.0000 347.6500 ;
      RECT 0.0000 347.2500 553.3800 347.5500 ;
      RECT 0.0000 345.5500 554.0000 347.2500 ;
      RECT 0.0000 345.2500 553.3800 345.5500 ;
      RECT 0.0000 344.3500 554.0000 345.2500 ;
      RECT 0.0000 344.0500 553.3800 344.3500 ;
      RECT 0.0000 341.9500 554.0000 344.0500 ;
      RECT 0.0000 341.6500 553.3800 341.9500 ;
      RECT 0.0000 340.7500 554.0000 341.6500 ;
      RECT 0.0000 340.4500 553.3800 340.7500 ;
      RECT 0.0000 338.3500 554.0000 340.4500 ;
      RECT 0.0000 338.0500 553.3800 338.3500 ;
      RECT 0.0000 337.1500 554.0000 338.0500 ;
      RECT 0.0000 336.8500 553.3800 337.1500 ;
      RECT 0.0000 334.7500 554.0000 336.8500 ;
      RECT 0.0000 334.4500 553.3800 334.7500 ;
      RECT 0.0000 333.5500 554.0000 334.4500 ;
      RECT 0.0000 333.2500 553.3800 333.5500 ;
      RECT 0.0000 329.9500 554.0000 333.2500 ;
      RECT 0.0000 329.6500 553.3800 329.9500 ;
      RECT 0.0000 329.5500 554.0000 329.6500 ;
      RECT 0.0000 329.2500 553.3800 329.5500 ;
      RECT 0.0000 322.7500 554.0000 329.2500 ;
      RECT 0.0000 322.4500 553.3800 322.7500 ;
      RECT 0.0000 308.3500 554.0000 322.4500 ;
      RECT 0.0000 308.0500 553.3800 308.3500 ;
      RECT 0.0000 307.9500 554.0000 308.0500 ;
      RECT 0.0000 307.6500 553.3800 307.9500 ;
      RECT 0.0000 304.9500 554.0000 307.6500 ;
      RECT 0.0000 304.6500 553.3800 304.9500 ;
      RECT 0.0000 302.3500 554.0000 304.6500 ;
      RECT 0.0000 302.0500 553.3800 302.3500 ;
      RECT 0.0000 295.1500 554.0000 302.0500 ;
      RECT 0.0000 294.8500 553.3800 295.1500 ;
      RECT 0.0000 294.3500 554.0000 294.8500 ;
      RECT 0.0000 294.0500 553.3800 294.3500 ;
      RECT 0.0000 293.9500 554.0000 294.0500 ;
      RECT 0.0000 293.6500 553.3800 293.9500 ;
      RECT 0.0000 293.5500 554.0000 293.6500 ;
      RECT 0.0000 293.2500 553.3800 293.5500 ;
      RECT 0.0000 283.1500 554.0000 293.2500 ;
      RECT 0.0000 282.8500 553.3800 283.1500 ;
      RECT 0.0000 280.7500 554.0000 282.8500 ;
      RECT 0.0000 280.4500 553.3800 280.7500 ;
      RECT 0.0000 275.9500 554.0000 280.4500 ;
      RECT 0.0000 275.6500 553.3800 275.9500 ;
      RECT 0.0000 273.5500 554.0000 275.6500 ;
      RECT 0.0000 273.2500 553.3800 273.5500 ;
      RECT 0.0000 273.1500 554.0000 273.2500 ;
      RECT 0.0000 272.8500 553.3800 273.1500 ;
      RECT 0.0000 272.3500 554.0000 272.8500 ;
      RECT 0.0000 272.0500 553.3800 272.3500 ;
      RECT 0.0000 271.9500 554.0000 272.0500 ;
      RECT 0.0000 271.6500 553.3800 271.9500 ;
      RECT 0.0000 269.9500 554.0000 271.6500 ;
      RECT 0.0000 269.6500 553.3800 269.9500 ;
      RECT 0.0000 268.7500 554.0000 269.6500 ;
      RECT 0.0000 268.4500 553.3800 268.7500 ;
      RECT 0.0000 266.3500 554.0000 268.4500 ;
      RECT 0.0000 266.0500 553.3800 266.3500 ;
      RECT 0.0000 265.1500 554.0000 266.0500 ;
      RECT 0.0000 264.8500 553.3800 265.1500 ;
      RECT 0.0000 261.9500 554.0000 264.8500 ;
      RECT 0.0000 261.6500 553.3800 261.9500 ;
      RECT 0.0000 261.5500 554.0000 261.6500 ;
      RECT 0.0000 261.2500 553.3800 261.5500 ;
      RECT 0.0000 261.1500 554.0000 261.2500 ;
      RECT 0.0000 260.8500 553.3800 261.1500 ;
      RECT 0.0000 257.9500 554.0000 260.8500 ;
      RECT 0.0000 257.6500 553.3800 257.9500 ;
      RECT 0.0000 255.5500 554.0000 257.6500 ;
      RECT 0.0000 255.2500 553.3800 255.5500 ;
      RECT 0.0000 251.9500 554.0000 255.2500 ;
      RECT 0.0000 251.6500 553.3800 251.9500 ;
      RECT 0.0000 250.7500 554.0000 251.6500 ;
      RECT 0.0000 250.4500 553.3800 250.7500 ;
      RECT 0.0000 250.3500 554.0000 250.4500 ;
      RECT 0.0000 250.0500 553.3800 250.3500 ;
      RECT 0.0000 248.3500 554.0000 250.0500 ;
      RECT 0.0000 248.0500 553.3800 248.3500 ;
      RECT 0.0000 243.5500 554.0000 248.0500 ;
      RECT 0.0000 243.2500 553.3800 243.5500 ;
      RECT 0.0000 241.1500 554.0000 243.2500 ;
      RECT 0.0000 240.8500 553.3800 241.1500 ;
      RECT 0.0000 240.7500 554.0000 240.8500 ;
      RECT 0.0000 240.4500 553.3800 240.7500 ;
      RECT 0.0000 239.9500 554.0000 240.4500 ;
      RECT 0.0000 239.6500 553.3800 239.9500 ;
      RECT 0.0000 237.5500 554.0000 239.6500 ;
      RECT 0.0000 237.2500 553.3800 237.5500 ;
      RECT 0.0000 232.7500 554.0000 237.2500 ;
      RECT 0.0000 232.4500 553.3800 232.7500 ;
      RECT 0.0000 227.9500 554.0000 232.4500 ;
      RECT 0.6200 227.6500 554.0000 227.9500 ;
      RECT 0.0000 225.5500 554.0000 227.6500 ;
      RECT 0.0000 225.2500 553.3800 225.5500 ;
      RECT 0.0000 225.1500 554.0000 225.2500 ;
      RECT 0.0000 224.8500 553.3800 225.1500 ;
      RECT 0.0000 223.1500 554.0000 224.8500 ;
      RECT 0.0000 222.8500 553.3800 223.1500 ;
      RECT 0.0000 220.5500 554.0000 222.8500 ;
      RECT 0.6200 220.2500 554.0000 220.5500 ;
      RECT 0.0000 219.9500 554.0000 220.2500 ;
      RECT 0.0000 219.6500 553.3800 219.9500 ;
      RECT 0.0000 219.5500 554.0000 219.6500 ;
      RECT 0.6200 219.2500 553.3800 219.5500 ;
      RECT 0.0000 219.1500 554.0000 219.2500 ;
      RECT 0.0000 218.8500 553.3800 219.1500 ;
      RECT 0.0000 218.3500 554.0000 218.8500 ;
      RECT 0.0000 218.0500 553.3800 218.3500 ;
      RECT 0.0000 217.9500 554.0000 218.0500 ;
      RECT 0.0000 217.6500 553.3800 217.9500 ;
      RECT 0.0000 217.3500 554.0000 217.6500 ;
      RECT 0.6200 217.0500 554.0000 217.3500 ;
      RECT 0.0000 216.7500 554.0000 217.0500 ;
      RECT 0.6200 216.4500 554.0000 216.7500 ;
      RECT 0.0000 216.1500 554.0000 216.4500 ;
      RECT 0.6200 215.9500 554.0000 216.1500 ;
      RECT 0.6200 215.8500 553.3800 215.9500 ;
      RECT 0.0000 215.7500 553.3800 215.8500 ;
      RECT 0.6200 215.6500 553.3800 215.7500 ;
      RECT 0.6200 215.5500 554.0000 215.6500 ;
      RECT 0.6200 215.4500 553.3800 215.5500 ;
      RECT 0.0000 215.3500 553.3800 215.4500 ;
      RECT 0.6200 215.2500 553.3800 215.3500 ;
      RECT 0.6200 215.0500 554.0000 215.2500 ;
      RECT 0.0000 213.3500 554.0000 215.0500 ;
      RECT 0.6200 213.0500 554.0000 213.3500 ;
      RECT 0.0000 211.3500 554.0000 213.0500 ;
      RECT 0.6200 211.0500 554.0000 211.3500 ;
      RECT 0.0000 210.7500 554.0000 211.0500 ;
      RECT 0.6200 210.4500 554.0000 210.7500 ;
      RECT 0.0000 210.3500 554.0000 210.4500 ;
      RECT 0.6200 210.0500 554.0000 210.3500 ;
      RECT 0.0000 209.9500 554.0000 210.0500 ;
      RECT 0.6200 209.6500 554.0000 209.9500 ;
      RECT 0.0000 209.5500 554.0000 209.6500 ;
      RECT 0.6200 209.2500 554.0000 209.5500 ;
      RECT 0.0000 208.5500 554.0000 209.2500 ;
      RECT 0.6200 208.2500 554.0000 208.5500 ;
      RECT 0.0000 205.9500 554.0000 208.2500 ;
      RECT 0.6200 205.6500 554.0000 205.9500 ;
      RECT 0.0000 205.3500 554.0000 205.6500 ;
      RECT 0.6200 205.0500 554.0000 205.3500 ;
      RECT 0.0000 204.3500 554.0000 205.0500 ;
      RECT 0.6200 204.0500 554.0000 204.3500 ;
      RECT 0.0000 203.5500 554.0000 204.0500 ;
      RECT 0.6200 203.2500 554.0000 203.5500 ;
      RECT 0.0000 201.3500 554.0000 203.2500 ;
      RECT 0.6200 201.0500 554.0000 201.3500 ;
      RECT 0.0000 198.9500 554.0000 201.0500 ;
      RECT 0.6200 198.6500 554.0000 198.9500 ;
      RECT 0.0000 198.5500 554.0000 198.6500 ;
      RECT 0.6200 198.2500 554.0000 198.5500 ;
      RECT 0.0000 198.1500 554.0000 198.2500 ;
      RECT 0.6200 197.8500 554.0000 198.1500 ;
      RECT 0.0000 196.1500 554.0000 197.8500 ;
      RECT 0.6200 195.8500 554.0000 196.1500 ;
      RECT 0.0000 195.5500 554.0000 195.8500 ;
      RECT 0.6200 195.2500 554.0000 195.5500 ;
      RECT 0.0000 195.1500 554.0000 195.2500 ;
      RECT 0.6200 194.8500 554.0000 195.1500 ;
      RECT 0.0000 194.3500 554.0000 194.8500 ;
      RECT 0.0000 194.0500 553.3800 194.3500 ;
      RECT 0.0000 193.7500 554.0000 194.0500 ;
      RECT 0.6200 193.4500 554.0000 193.7500 ;
      RECT 0.0000 193.1500 554.0000 193.4500 ;
      RECT 0.0000 192.8500 553.3800 193.1500 ;
      RECT 0.0000 192.7500 554.0000 192.8500 ;
      RECT 0.0000 192.4500 553.3800 192.7500 ;
      RECT 0.0000 191.7500 554.0000 192.4500 ;
      RECT 0.6200 191.4500 554.0000 191.7500 ;
      RECT 0.0000 186.7500 554.0000 191.4500 ;
      RECT 0.6200 186.4500 554.0000 186.7500 ;
      RECT 0.0000 185.9500 554.0000 186.4500 ;
      RECT 0.0000 185.6500 553.3800 185.9500 ;
      RECT 0.0000 172.7500 554.0000 185.6500 ;
      RECT 0.0000 172.4500 553.3800 172.7500 ;
      RECT 0.0000 146.3500 554.0000 172.4500 ;
      RECT 0.0000 146.0500 553.3800 146.3500 ;
      RECT 0.0000 140.3500 554.0000 146.0500 ;
      RECT 0.0000 140.0500 553.3800 140.3500 ;
      RECT 0.0000 134.3500 554.0000 140.0500 ;
      RECT 0.6200 134.0500 554.0000 134.3500 ;
      RECT 0.0000 131.5500 554.0000 134.0500 ;
      RECT 0.6200 131.2500 554.0000 131.5500 ;
      RECT 0.0000 128.3500 554.0000 131.2500 ;
      RECT 0.0000 128.0500 553.3800 128.3500 ;
      RECT 0.0000 120.5500 554.0000 128.0500 ;
      RECT 0.6200 120.2500 554.0000 120.5500 ;
      RECT 0.0000 118.1500 554.0000 120.2500 ;
      RECT 0.6200 117.8500 554.0000 118.1500 ;
      RECT 0.0000 113.9500 554.0000 117.8500 ;
      RECT 0.0000 113.6500 553.3800 113.9500 ;
      RECT 0.0000 107.9500 554.0000 113.6500 ;
      RECT 0.0000 107.6500 553.3800 107.9500 ;
      RECT 0.0000 96.3500 554.0000 107.6500 ;
      RECT 0.6200 96.0500 554.0000 96.3500 ;
      RECT 0.0000 92.1500 554.0000 96.0500 ;
      RECT 0.6200 91.8500 554.0000 92.1500 ;
      RECT 0.0000 91.7500 554.0000 91.8500 ;
      RECT 0.6200 91.4500 554.0000 91.7500 ;
      RECT 0.0000 86.3500 554.0000 91.4500 ;
      RECT 0.6200 86.0500 554.0000 86.3500 ;
      RECT 0.0000 76.3500 554.0000 86.0500 ;
      RECT 0.6200 76.0500 554.0000 76.3500 ;
      RECT 0.0000 73.9500 554.0000 76.0500 ;
      RECT 0.6200 73.6500 554.0000 73.9500 ;
      RECT 0.0000 72.9500 554.0000 73.6500 ;
      RECT 0.6200 72.6500 554.0000 72.9500 ;
      RECT 0.0000 72.3500 554.0000 72.6500 ;
      RECT 0.6200 72.0500 554.0000 72.3500 ;
      RECT 0.0000 71.9500 554.0000 72.0500 ;
      RECT 0.6200 71.6500 554.0000 71.9500 ;
      RECT 0.0000 71.5500 554.0000 71.6500 ;
      RECT 0.6200 71.2500 554.0000 71.5500 ;
      RECT 0.0000 57.3500 554.0000 71.2500 ;
      RECT 0.6200 57.0500 554.0000 57.3500 ;
      RECT 0.0000 0.0000 554.0000 57.0500 ;
    LAYER M4 ;
      RECT 519.2500 550.5000 535.7500 551.0000 ;
      RECT 0.0000 550.5000 510.5500 551.0000 ;
      RECT 536.0500 550.3800 554.0000 551.0000 ;
      RECT 527.4900 550.3800 535.7500 550.5000 ;
      RECT 519.2500 550.3800 524.4900 550.5000 ;
      RECT 510.8500 550.3800 518.9500 551.0000 ;
      RECT 499.4350 550.3800 510.5500 550.5000 ;
      RECT 527.4900 545.5000 554.0000 550.3800 ;
      RECT 499.4350 545.5000 524.4900 550.3800 ;
      RECT 471.3800 545.5000 496.4350 550.5000 ;
      RECT 443.3250 545.5000 468.3800 550.5000 ;
      RECT 415.2700 545.5000 440.3250 550.5000 ;
      RECT 387.2150 545.5000 412.2700 550.5000 ;
      RECT 359.1600 545.5000 384.2150 550.5000 ;
      RECT 331.1050 545.5000 356.1600 550.5000 ;
      RECT 303.0500 545.5000 328.1050 550.5000 ;
      RECT 274.9950 545.5000 300.0500 550.5000 ;
      RECT 246.9400 545.5000 271.9950 550.5000 ;
      RECT 218.8850 545.5000 243.9400 550.5000 ;
      RECT 190.8300 545.5000 215.8850 550.5000 ;
      RECT 162.7750 545.5000 187.8300 550.5000 ;
      RECT 134.7200 545.5000 159.7750 550.5000 ;
      RECT 106.6650 545.5000 131.7200 550.5000 ;
      RECT 78.6100 545.5000 103.6650 550.5000 ;
      RECT 50.5550 545.5000 75.6100 550.5000 ;
      RECT 22.5000 545.5000 47.5550 550.5000 ;
      RECT 535.4900 5.5000 554.0000 545.5000 ;
      RECT 527.4900 5.5000 532.4900 545.5000 ;
      RECT 507.4350 5.5000 524.4900 545.5000 ;
      RECT 499.4350 5.5000 504.4350 545.5000 ;
      RECT 479.3800 5.5000 496.4350 545.5000 ;
      RECT 471.3800 5.5000 476.3800 545.5000 ;
      RECT 451.3250 5.5000 468.3800 545.5000 ;
      RECT 443.3250 5.5000 448.3250 545.5000 ;
      RECT 423.2700 5.5000 440.3250 545.5000 ;
      RECT 415.2700 5.5000 420.2700 545.5000 ;
      RECT 395.2150 5.5000 412.2700 545.5000 ;
      RECT 387.2150 5.5000 392.2150 545.5000 ;
      RECT 367.1600 5.5000 384.2150 545.5000 ;
      RECT 359.1600 5.5000 364.1600 545.5000 ;
      RECT 339.1050 5.5000 356.1600 545.5000 ;
      RECT 331.1050 5.5000 336.1050 545.5000 ;
      RECT 311.0500 5.5000 328.1050 545.5000 ;
      RECT 303.0500 5.5000 308.0500 545.5000 ;
      RECT 282.9950 5.5000 300.0500 545.5000 ;
      RECT 274.9950 5.5000 279.9950 545.5000 ;
      RECT 254.9400 5.5000 271.9950 545.5000 ;
      RECT 246.9400 5.5000 251.9400 545.5000 ;
      RECT 226.8850 5.5000 243.9400 545.5000 ;
      RECT 218.8850 5.5000 223.8850 545.5000 ;
      RECT 198.8300 5.5000 215.8850 545.5000 ;
      RECT 190.8300 5.5000 195.8300 545.5000 ;
      RECT 170.7750 5.5000 187.8300 545.5000 ;
      RECT 162.7750 5.5000 167.7750 545.5000 ;
      RECT 142.7200 5.5000 159.7750 545.5000 ;
      RECT 134.7200 5.5000 139.7200 545.5000 ;
      RECT 114.6650 5.5000 131.7200 545.5000 ;
      RECT 106.6650 5.5000 111.6650 545.5000 ;
      RECT 86.6100 5.5000 103.6650 545.5000 ;
      RECT 78.6100 5.5000 83.6100 545.5000 ;
      RECT 58.5550 5.5000 75.6100 545.5000 ;
      RECT 50.5550 5.5000 55.5550 545.5000 ;
      RECT 30.5000 5.5000 47.5550 545.5000 ;
      RECT 22.5000 5.5000 27.5000 545.5000 ;
      RECT 471.3800 0.6200 496.4350 5.5000 ;
      RECT 162.7750 0.6200 187.8300 5.5000 ;
      RECT 527.4900 0.5000 554.0000 5.5000 ;
      RECT 499.4350 0.5000 524.4900 5.5000 ;
      RECT 485.8500 0.5000 496.4350 0.6200 ;
      RECT 471.3800 0.5000 477.1500 0.6200 ;
      RECT 443.3250 0.5000 468.3800 5.5000 ;
      RECT 415.2700 0.5000 440.3250 5.5000 ;
      RECT 387.2150 0.5000 412.2700 5.5000 ;
      RECT 359.1600 0.5000 384.2150 5.5000 ;
      RECT 331.1050 0.5000 356.1600 5.5000 ;
      RECT 303.0500 0.5000 328.1050 5.5000 ;
      RECT 274.9950 0.5000 300.0500 5.5000 ;
      RECT 246.9400 0.5000 271.9950 5.5000 ;
      RECT 218.8850 0.5000 243.9400 5.5000 ;
      RECT 190.8300 0.5000 215.8850 5.5000 ;
      RECT 165.0500 0.5000 187.8300 0.6200 ;
      RECT 162.7750 0.5000 164.7500 0.6200 ;
      RECT 134.7200 0.5000 159.7750 5.5000 ;
      RECT 106.6650 0.5000 131.7200 5.5000 ;
      RECT 78.6100 0.5000 103.6650 5.5000 ;
      RECT 50.5550 0.5000 75.6100 5.5000 ;
      RECT 22.5000 0.5000 47.5550 5.5000 ;
      RECT 0.0000 0.5000 19.5000 550.5000 ;
      RECT 485.8500 0.0000 554.0000 0.5000 ;
      RECT 477.4500 0.0000 485.5500 0.6200 ;
      RECT 165.0500 0.0000 477.1500 0.5000 ;
      RECT 0.0000 0.0000 164.7500 0.5000 ;
  END
END fullchip

END LIBRARY
